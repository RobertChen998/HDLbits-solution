`timescale 1ns/10ps

module tb();

    reg               clk;
    reg               i_rst_n;
    reg               i_inhibit;
    reg               i_valid;
    reg      [ 9-1:0] i_q;	// Need to handle at last, we now use the difference and pipeline to the last stage...
    reg      [ 9-1:0] zero_vector;

    reg      [ 8-1:0] i_im1;
    reg      [ 8-1:0] i_im2;
    reg      [ 8-1:0] i_im3;
    reg      [ 8-1:0] i_im4;
    reg      [ 8-1:0] i_im5;
    reg      [ 8-1:0] i_im6;
    reg      [ 8-1:0] i_im7;
    reg      [ 8-1:0] i_im8;
    reg      [ 8-1:0] i_im9;

    reg      [ 4-1:0] i_ker1;
    reg      [ 4-1:0] i_ker2;
    reg      [ 4-1:0] i_ker3;
    reg      [ 4-1:0] i_ker4;
    reg      [ 4-1:0] i_ker5;
    reg      [ 4-1:0] i_ker6;
    reg      [ 4-1:0] i_ker7;
    reg      [ 4-1:0] i_ker8;
    reg      [ 4-1:0] i_ker9;

    wire             o_valid;
    wire     [15:0]   o_conv;

    initial begin
        $dumpfile("mac.fsdb");
        $dumpvars;
        clk = 1'b0;
        i_rst_n = 1'b1;
        i_valid = 1'b0;
        i_inhibit = 1'b0;

        // i_im1 = 8'b00110111;
        // i_im2 = 8'b00110000;
        // i_im3 = 8'b00111000;
        // i_im4 = 8'b00111100;
        // i_im5 = 8'b00110101;
        // i_im6 = 8'b00110111;
        // i_im7 = 8'b00100111;
        // i_im8 = 8'b00111010;
        // i_im9 = 8'b00110110;

        // 1-1
        i_im1 = 8'h3C;
        i_im2 = 8'h37;
        i_im3 = 8'hB6;
        i_im4 = 8'h35;
        i_im5 = 8'h36;
        i_im6 = 8'hBB;
        i_im7 = 8'h38;
        i_im8 = 8'hA6;
        i_im9 = 8'hB2;


// =============  i_ker  =================== //
        // i_ker1 = 4'b0010;
        // i_ker2 = 4'b0001;
        // i_ker3 = 4'b1010;
        // i_ker4 = 4'b0110;
        // i_ker5 = 4'b1001;
        // i_ker6 = 4'b0110;
        // i_ker7 = 4'b1011;
        // i_ker8 = 4'b0001;
        // i_ker9 = 4'b0101;
        
        i_ker1 = 4'hB;
        i_ker2 = 4'hC;
        i_ker3 = 4'hC;
        i_ker4 = 4'hD;
        i_ker5 = 4'hD;
        i_ker6 = 4'hE;
        i_ker7 = 4'h3;
        i_ker8 = 4'h5;
        i_ker9 = 4'h5;

        #1 i_rst_n = 1'b0;
        #5 i_rst_n = 1'b1;
        #20 i_valid = 1'b1;

        #10 //1-2
        i_im1 = 8'h37;
        i_im2 = 8'hB6;
        i_im3 = 8'hA8;
        i_im4 = 8'h36;
        i_im5 = 8'hBB;
        i_im6 = 8'h39;
        i_im7 = 8'hA6;
        i_im8 = 8'hB2;
        i_im9 = 8'hAF;

        #10 //1-3
        i_im1 = 8'hB6;
        i_im2 = 8'hA8;
        i_im3 = 8'h3C;
        i_im4 = 8'hBB;
        i_im5 = 8'h39;
        i_im6 = 8'h31;
        i_im7 = 8'hB2;
        i_im8 = 8'hAF;
        i_im9 = 8'hB8;
        #10 //1-4
        i_im1 = 8'hA8;
        i_im2 = 8'h3C;
        i_im3 = 8'h33;
        i_im4 = 8'h39;
        i_im5 = 8'h31;
        i_im6 = 8'hB6;
        i_im7 = 8'hAF;
        i_im8 = 8'hB8;
        i_im9 = 8'hB3;
        #10 //1-5
        i_im1 = 8'h3C;
        i_im2 = 8'h33;
        i_im3 = 8'h3C;
        i_im4 = 8'h31;
        i_im5 = 8'hB6;
        i_im6 = 8'hBC;
        i_im7 = 8'hB8;
        i_im8 = 8'hB3;
        i_im9 = 8'hB2;
        #10 //1-6
        i_im1 = 8'h33;
        i_im2 = 8'h3C;
        i_im3 = 8'hB6;
        i_im4 = 8'hB6;
        i_im5 = 8'hBC;
        i_im6 = 8'h36;
        i_im7 = 8'hB3;
        i_im8 = 8'hB2;
        i_im9 = 8'hAF;
        #10 //1-7
        i_im1 = 8'h3C;
        i_im2 = 8'hB6;
        i_im3 = 8'hB6;
        i_im4 = 8'hBC;
        i_im5 = 8'h36;
        i_im6 = 8'h3A;
        i_im7 = 8'hB2;
        i_im8 = 8'hAF;
        i_im9 = 8'h38;
        #10 //1-8
        i_im1 = 8'hB6;
        i_im2 = 8'hB6;
        i_im3 = 8'h3A;
        i_im4 = 8'h36;
        i_im5 = 8'h3A;
        i_im6 = 8'h3B;
        i_im7 = 8'hAF;
        i_im8 = 8'h38;
        i_im9 = 8'h3A;
        #10 //1-9
        i_im1 = 8'hB6;
        i_im2 = 8'h3A;
        i_im3 = 8'hB6;
        i_im4 = 8'h3A;
        i_im5 = 8'h3B;
        i_im6 = 8'h37;
        i_im7 = 8'h38;
        i_im8 = 8'h3A;
        i_im9 = 8'hB4;
        #10 //1-10
        i_im1 = 8'h3A;
        i_im2 = 8'hB6;
        i_im3 = 8'hBB;
        i_im4 = 8'h3B;
        i_im5 = 8'h37;
        i_im6 = 8'hB6;
        i_im7 = 8'h3A;
        i_im8 = 8'hB4;
        i_im9 = 8'hB8;
        #10 //1-11
        i_im1 = 8'hB6;
        i_im2 = 8'hBB;
        i_im3 = 8'hB9;
        i_im4 = 8'h37;
        i_im5 = 8'hB6;
        i_im6 = 8'hB8;
        i_im7 = 8'hB4;
        i_im8 = 8'hB8;
        i_im9 = 8'h3A;
        #10 //1-12
        i_im1 = 8'hBB;
        i_im2 = 8'hB9;
        i_im3 = 8'h35;
        i_im4 = 8'hB6;
        i_im5 = 8'hB8;
        i_im6 = 8'hBB;
        i_im7 = 8'hB8;
        i_im8 = 8'h3A;
        i_im9 = 8'hBA;
        #10 //1-13
        i_im1 = 8'hB9;
        i_im2 = 8'h35;
        i_im3 = 8'hBC;
        i_im4 = 8'hB8;
        i_im5 = 8'hBB;
        i_im6 = 8'h33;
        i_im7 = 8'h3A;
        i_im8 = 8'hBA;
        i_im9 = 8'h3B;
        #10 //1-14
        i_im1 = 8'h35;
        i_im2 = 8'hBC;
        i_im3 = 8'hB2;
        i_im4 = 8'hBB;
        i_im5 = 8'h33;
        i_im6 = 8'hBA;
        i_im7 = 8'hBA;
        i_im8 = 8'h3B;
        i_im9 = 8'hBA;
        #10 //1-15
        i_im1 = 8'hBC;
        i_im2 = 8'hB2;
        i_im3 = 8'h38;
        i_im4 = 8'h33;
        i_im5 = 8'hBA;
        i_im6 = 8'hBB;
        i_im7 = 8'h3B;
        i_im8 = 8'hBA;
        i_im9 = 8'hB9;
        #10 //1-16
        i_im1 = 8'hB2;
        i_im2 = 8'h38;
        i_im3 = 8'h38;
        i_im4 = 8'hBA;
        i_im5 = 8'hBB;
        i_im6 = 8'h34;
        i_im7 = 8'hBA;
        i_im8 = 8'hB9;
        i_im9 = 8'h27;
        #10 //1-17
        i_im1 = 8'h38;
        i_im2 = 8'h38;
        i_im3 = 8'hB7;
        i_im4 = 8'hBB;
        i_im5 = 8'h34;
        i_im6 = 8'hA9;
        i_im7 = 8'hB9;
        i_im8 = 8'h27;
        i_im9 = 8'h3B;
        #10 //1-18
        i_im1 = 8'h38;
        i_im2 = 8'hB7;
        i_im3 = 8'hB9;
        i_im4 = 8'h34;
        i_im5 = 8'hA9;
        i_im6 = 8'h36;
        i_im7 = 8'h27;
        i_im8 = 8'h3B;
        i_im9 = 8'h39;
        #10 //1-19
        i_im1 = 8'hB7;
        i_im2 = 8'hB9;
        i_im3 = 8'h3B;
        i_im4 = 8'hA9;
        i_im5 = 8'h36;
        i_im6 = 8'h37;
        i_im7 = 8'h3B;
        i_im8 = 8'h39;
        i_im9 = 8'h3B;
        #10 //1-20
        i_im1 = 8'hB9;
        i_im2 = 8'h3B;
        i_im3 = 8'h39;
        i_im4 = 8'h36;
        i_im5 = 8'h37;
        i_im6 = 8'hB5;
        i_im7 = 8'h39;
        i_im8 = 8'h3B;
        i_im9 = 8'hB8;
        #10 //1-21
        i_im1 = 8'h3B;
        i_im2 = 8'h39;
        i_im3 = 8'hB9;
        i_im4 = 8'h37;
        i_im5 = 8'hB5;
        i_im6 = 8'hB9;
        i_im7 = 8'h3B;
        i_im8 = 8'hB8;
        i_im9 = 8'h3B;
        #10 //1-22
        i_im1 = 8'h39;
        i_im2 = 8'hB9;
        i_im3 = 8'hB7;
        i_im4 = 8'hB5;
        i_im5 = 8'hB9;
        i_im6 = 8'h2D;
        i_im7 = 8'hB8;
        i_im8 = 8'h3B;
        i_im9 = 8'hAF;
        #10 //1-23
        i_im1 = 8'hB9;
        i_im2 = 8'hB7;
        i_im3 = 8'hB1;
        i_im4 = 8'hB9;
        i_im5 = 8'h2D;
        i_im6 = 8'hA2;
        i_im7 = 8'h3B;
        i_im8 = 8'hAF;
        i_im9 = 8'hBA;
        #10 //1-24
        i_im1 = 8'hB7;
        i_im2 = 8'hB1;
        i_im3 = 8'hBC;
        i_im4 = 8'h2D;
        i_im5 = 8'hA2;
        i_im6 = 8'hBC;
        i_im7 = 8'hAF;
        i_im8 = 8'hBA;
        i_im9 = 8'h38;
        #10 //1-25
        i_im1 = 8'hB1;
        i_im2 = 8'hBC;
        i_im3 = 8'hB9;
        i_im4 = 8'hA2;
        i_im5 = 8'hBC;
        i_im6 = 8'h29;
        i_im7 = 8'hBA;
        i_im8 = 8'h38;
        i_im9 = 8'h2B;
        #10 //1-26
        i_im1 = 8'hBC;
        i_im2 = 8'hB9;
        i_im3 = 8'hB8;
        i_im4 = 8'hBC;
        i_im5 = 8'h29;
        i_im6 = 8'h39;
        i_im7 = 8'h38;
        i_im8 = 8'h2B;
        i_im9 = 8'h34;
        #10 //2-1
        i_im1 = 8'h35;
        i_im2 = 8'h36;
        i_im3 = 8'hBB;
        i_im4 = 8'h38;
        i_im5 = 8'hA6;
        i_im6 = 8'hB2;
        i_im7 = 8'hB4;
        i_im8 = 8'hB5;
        i_im9 = 8'hB9;
        #10 //2-2
        i_im1 = 8'h36;
        i_im2 = 8'hBB;
        i_im3 = 8'h39;
        i_im4 = 8'hA6;
        i_im5 = 8'hB2;
        i_im6 = 8'hAF;
        i_im7 = 8'hB5;
        i_im8 = 8'hB9;
        i_im9 = 8'hB7;
        #10 //2-3
        i_im1 = 8'hBB;
        i_im2 = 8'h39;
        i_im3 = 8'h31;
        i_im4 = 8'hB2;
        i_im5 = 8'hAF;
        i_im6 = 8'hB8;
        i_im7 = 8'hB9;
        i_im8 = 8'hB7;
        i_im9 = 8'hB5;
        #10 //2-4
        i_im1 = 8'h39;
        i_im2 = 8'h31;
        i_im3 = 8'hB6;
        i_im4 = 8'hAF;
        i_im5 = 8'hB8;
        i_im6 = 8'hB3;
        i_im7 = 8'hB7;
        i_im8 = 8'hB5;
        i_im9 = 8'hB7;
        #10 //2-5
        i_im1 = 8'h31;
        i_im2 = 8'hB6;
        i_im3 = 8'hBC;
        i_im4 = 8'hB8;
        i_im5 = 8'hB3;
        i_im6 = 8'hB2;
        i_im7 = 8'hB5;
        i_im8 = 8'hB7;
        i_im9 = 8'hB4;
        #10 //2-6
        i_im1 = 8'hB6;
        i_im2 = 8'hBC;
        i_im3 = 8'h36;
        i_im4 = 8'hB3;
        i_im5 = 8'hB2;
        i_im6 = 8'hAF;
        i_im7 = 8'hB7;
        i_im8 = 8'hB4;
        i_im9 = 8'h3A;
        #10 //2-7
        i_im1 = 8'hBC;
        i_im2 = 8'h36;
        i_im3 = 8'h3A;
        i_im4 = 8'hB2;
        i_im5 = 8'hAF;
        i_im6 = 8'h38;
        i_im7 = 8'hB4;
        i_im8 = 8'h3A;
        i_im9 = 8'hBB;
        #10 //2-8
        i_im1 = 8'h36;
        i_im2 = 8'h3A;
        i_im3 = 8'h3B;
        i_im4 = 8'hAF;
        i_im5 = 8'h38;
        i_im6 = 8'h3A;
        i_im7 = 8'h3A;
        i_im8 = 8'hBB;
        i_im9 = 8'hB8;
        #10 //2-9
        i_im1 = 8'h3A;
        i_im2 = 8'h3B;
        i_im3 = 8'h37;
        i_im4 = 8'h38;
        i_im5 = 8'h3A;
        i_im6 = 8'hB4;
        i_im7 = 8'hBB;
        i_im8 = 8'hB8;
        i_im9 = 8'hB1;
        #10 //2-10
        i_im1 = 8'h3B;
        i_im2 = 8'h37;
        i_im3 = 8'hB6;
        i_im4 = 8'h3A;
        i_im5 = 8'hB4;
        i_im6 = 8'hB8;
        i_im7 = 8'hB8;
        i_im8 = 8'hB1;
        i_im9 = 8'hB2;
        #10 //2-11
        i_im1 = 8'h37;
        i_im2 = 8'hB6;
        i_im3 = 8'hB8;
        i_im4 = 8'hB4;
        i_im5 = 8'hB8;
        i_im6 = 8'h3A;
        i_im7 = 8'hB1;
        i_im8 = 8'hB2;
        i_im9 = 8'hB2;
        #10 //2-12
        i_im1 = 8'hB6;
        i_im2 = 8'hB8;
        i_im3 = 8'hBB;
        i_im4 = 8'hB8;
        i_im5 = 8'h3A;
        i_im6 = 8'hBA;
        i_im7 = 8'hB2;
        i_im8 = 8'hB2;
        i_im9 = 8'hB8;
        #10 //2-13
        i_im1 = 8'hB8;
        i_im2 = 8'hBB;
        i_im3 = 8'h33;
        i_im4 = 8'h3A;
        i_im5 = 8'hBA;
        i_im6 = 8'h3B;
        i_im7 = 8'hB2;
        i_im8 = 8'hB8;
        i_im9 = 8'h39;
        #10 //2-14
        i_im1 = 8'hBB;
        i_im2 = 8'h33;
        i_im3 = 8'hBA;
        i_im4 = 8'hBA;
        i_im5 = 8'h3B;
        i_im6 = 8'hBA;
        i_im7 = 8'hB8;
        i_im8 = 8'h39;
        i_im9 = 8'h39;
        #10 //2-15
        i_im1 = 8'h33;
        i_im2 = 8'hBA;
        i_im3 = 8'hBB;
        i_im4 = 8'h3B;
        i_im5 = 8'hBA;
        i_im6 = 8'hB9;
        i_im7 = 8'h39;
        i_im8 = 8'h39;
        i_im9 = 8'hBB;
        #10 //2-16
        i_im1 = 8'hBA;
        i_im2 = 8'hBB;
        i_im3 = 8'h34;
        i_im4 = 8'hBA;
        i_im5 = 8'hB9;
        i_im6 = 8'h27;
        i_im7 = 8'h39;
        i_im8 = 8'hBB;
        i_im9 = 8'hB7;
        #10 //2-17
        i_im1 = 8'hBB;
        i_im2 = 8'h34;
        i_im3 = 8'hA9;
        i_im4 = 8'hB9;
        i_im5 = 8'h27;
        i_im6 = 8'h3B;
        i_im7 = 8'hBB;
        i_im8 = 8'hB7;
        i_im9 = 8'h35;
        #10 //2-18
        i_im1 = 8'h34;
        i_im2 = 8'hA9;
        i_im3 = 8'h36;
        i_im4 = 8'h27;
        i_im5 = 8'h3B;
        i_im6 = 8'h39;
        i_im7 = 8'hB7;
        i_im8 = 8'h35;
        i_im9 = 8'h35;
        #10 //2-19
        i_im1 = 8'hA9;
        i_im2 = 8'h36;
        i_im3 = 8'h37;
        i_im4 = 8'h3B;
        i_im5 = 8'h39;
        i_im6 = 8'h3B;
        i_im7 = 8'h35;
        i_im8 = 8'h35;
        i_im9 = 8'hBB;
        #10 //2-20
        i_im1 = 8'h36;
        i_im2 = 8'h37;
        i_im3 = 8'hB5;
        i_im4 = 8'h39;
        i_im5 = 8'h3B;
        i_im6 = 8'hB8;
        i_im7 = 8'h35;
        i_im8 = 8'hBB;
        i_im9 = 8'h20;
        #10 //2-21
        i_im1 = 8'h37;
        i_im2 = 8'hB5;
        i_im3 = 8'hB9;
        i_im4 = 8'h3B;
        i_im5 = 8'hB8;
        i_im6 = 8'h3B;
        i_im7 = 8'hBB;
        i_im8 = 8'h20;
        i_im9 = 8'h35;
        #10 //2-22
        i_im1 = 8'hB5;
        i_im2 = 8'hB9;
        i_im3 = 8'h2D;
        i_im4 = 8'hB8;
        i_im5 = 8'h3B;
        i_im6 = 8'hAF;
        i_im7 = 8'h20;
        i_im8 = 8'h35;
        i_im9 = 8'hB9;
        #10 //2-23
        i_im1 = 8'hB9;
        i_im2 = 8'h2D;
        i_im3 = 8'hA2;
        i_im4 = 8'h3B;
        i_im5 = 8'hAF;
        i_im6 = 8'hBA;
        i_im7 = 8'h35;
        i_im8 = 8'hB9;
        i_im9 = 8'h39;
        #10 //2-24
        i_im1 = 8'h2D;
        i_im2 = 8'hA2;
        i_im3 = 8'hBC;
        i_im4 = 8'hAF;
        i_im5 = 8'hBA;
        i_im6 = 8'h38;
        i_im7 = 8'hB9;
        i_im8 = 8'h39;
        i_im9 = 8'hB1;
        #10 //2-25
        i_im1 = 8'hA2;
        i_im2 = 8'hBC;
        i_im3 = 8'h29;
        i_im4 = 8'hBA;
        i_im5 = 8'h38;
        i_im6 = 8'h2B;
        i_im7 = 8'h39;
        i_im8 = 8'hB1;
        i_im9 = 8'hBB;
        #10 //2-26
        i_im1 = 8'hBC;
        i_im2 = 8'h29;
        i_im3 = 8'h39;
        i_im4 = 8'h38;
        i_im5 = 8'h2B;
        i_im6 = 8'h34;
        i_im7 = 8'hB1;
        i_im8 = 8'hBB;
        i_im9 = 8'h30;
        #10 //3-1
        i_im1 = 8'h38;
        i_im2 = 8'hA6;
        i_im3 = 8'hB2;
        i_im4 = 8'hB4;
        i_im5 = 8'hB5;
        i_im6 = 8'hB9;
        i_im7 = 8'hBB;
        i_im8 = 8'h3A;
        i_im9 = 8'h39;
        #10 //3-2
        i_im1 = 8'hA6;
        i_im2 = 8'hB2;
        i_im3 = 8'hAF;
        i_im4 = 8'hB5;
        i_im5 = 8'hB9;
        i_im6 = 8'hB7;
        i_im7 = 8'h3A;
        i_im8 = 8'h39;
        i_im9 = 8'h37;
        #10 //3-3
        i_im1 = 8'hB2;
        i_im2 = 8'hAF;
        i_im3 = 8'hB8;
        i_im4 = 8'hB9;
        i_im5 = 8'hB7;
        i_im6 = 8'hB5;
        i_im7 = 8'h39;
        i_im8 = 8'h37;
        i_im9 = 8'hB7;
        #10 //3-4
        i_im1 = 8'hAF;
        i_im2 = 8'hB8;
        i_im3 = 8'hB3;
        i_im4 = 8'hB7;
        i_im5 = 8'hB5;
        i_im6 = 8'hB7;
        i_im7 = 8'h37;
        i_im8 = 8'hB7;
        i_im9 = 8'h3A;
        #10 //3-5
        i_im1 = 8'hB8;
        i_im2 = 8'hB3;
        i_im3 = 8'hB2;
        i_im4 = 8'hB5;
        i_im5 = 8'hB7;
        i_im6 = 8'hB4;
        i_im7 = 8'hB7;
        i_im8 = 8'h3A;
        i_im9 = 8'h20;
        #10 //3-6
        i_im1 = 8'hB3;
        i_im2 = 8'hB2;
        i_im3 = 8'hAF;
        i_im4 = 8'hB7;
        i_im5 = 8'hB4;
        i_im6 = 8'h3A;
        i_im7 = 8'h3A;
        i_im8 = 8'h20;
        i_im9 = 8'hBB;
        #10 //3-7
        i_im1 = 8'hB2;
        i_im2 = 8'hAF;
        i_im3 = 8'h38;
        i_im4 = 8'hB4;
        i_im5 = 8'h3A;
        i_im6 = 8'hBB;
        i_im7 = 8'h20;
        i_im8 = 8'hBB;
        i_im9 = 8'hB9;
        #10 //3-8
        i_im1 = 8'hAF;
        i_im2 = 8'h38;
        i_im3 = 8'h3A;
        i_im4 = 8'h3A;
        i_im5 = 8'hBB;
        i_im6 = 8'hB8;
        i_im7 = 8'hBB;
        i_im8 = 8'hB9;
        i_im9 = 8'h29;
        #10 //3-9
        i_im1 = 8'h38;
        i_im2 = 8'h3A;
        i_im3 = 8'hB4;
        i_im4 = 8'hBB;
        i_im5 = 8'hB8;
        i_im6 = 8'hB1;
        i_im7 = 8'hB9;
        i_im8 = 8'h29;
        i_im9 = 8'hB8;
        #10 //3-10
        i_im1 = 8'h3A;
        i_im2 = 8'hB4;
        i_im3 = 8'hB8;
        i_im4 = 8'hB8;
        i_im5 = 8'hB1;
        i_im6 = 8'hB2;
        i_im7 = 8'h29;
        i_im8 = 8'hB8;
        i_im9 = 8'hB1;
        #10 //3-11
        i_im1 = 8'hB4;
        i_im2 = 8'hB8;
        i_im3 = 8'h3A;
        i_im4 = 8'hB1;
        i_im5 = 8'hB2;
        i_im6 = 8'hB2;
        i_im7 = 8'hB8;
        i_im8 = 8'hB1;
        i_im9 = 8'hA5;
        #10 //3-12
        i_im1 = 8'hB8;
        i_im2 = 8'h3A;
        i_im3 = 8'hBA;
        i_im4 = 8'hB2;
        i_im5 = 8'hB2;
        i_im6 = 8'hB8;
        i_im7 = 8'hB1;
        i_im8 = 8'hA5;
        i_im9 = 8'hBA;
        #10 //3-13
        i_im1 = 8'h3A;
        i_im2 = 8'hBA;
        i_im3 = 8'h3B;
        i_im4 = 8'hB2;
        i_im5 = 8'hB8;
        i_im6 = 8'h39;
        i_im7 = 8'hA5;
        i_im8 = 8'hBA;
        i_im9 = 8'hBA;
        #10 //3-14
        i_im1 = 8'hBA;
        i_im2 = 8'h3B;
        i_im3 = 8'hBA;
        i_im4 = 8'hB8;
        i_im5 = 8'h39;
        i_im6 = 8'h39;
        i_im7 = 8'hBA;
        i_im8 = 8'hBA;
        i_im9 = 8'h30;
        #10 //3-15
        i_im1 = 8'h3B;
        i_im2 = 8'hBA;
        i_im3 = 8'hB9;
        i_im4 = 8'h39;
        i_im5 = 8'h39;
        i_im6 = 8'hBB;
        i_im7 = 8'hBA;
        i_im8 = 8'h30;
        i_im9 = 8'h36;
        #10 //3-16
        i_im1 = 8'hBA;
        i_im2 = 8'hB9;
        i_im3 = 8'h27;
        i_im4 = 8'h39;
        i_im5 = 8'hBB;
        i_im6 = 8'hB7;
        i_im7 = 8'h30;
        i_im8 = 8'h36;
        i_im9 = 8'hB9;
        #10 //3-17
        i_im1 = 8'hB9;
        i_im2 = 8'h27;
        i_im3 = 8'h3B;
        i_im4 = 8'hBB;
        i_im5 = 8'hB7;
        i_im6 = 8'h35;
        i_im7 = 8'h36;
        i_im8 = 8'hB9;
        i_im9 = 8'hA8;
        #10 //3-18
        i_im1 = 8'h27;
        i_im2 = 8'h3B;
        i_im3 = 8'h39;
        i_im4 = 8'hB7;
        i_im5 = 8'h35;
        i_im6 = 8'h35;
        i_im7 = 8'hB9;
        i_im8 = 8'hA8;
        i_im9 = 8'hB8;
        #10 //3-19
        i_im1 = 8'h3B;
        i_im2 = 8'h39;
        i_im3 = 8'h3B;
        i_im4 = 8'h35;
        i_im5 = 8'h35;
        i_im6 = 8'hBB;
        i_im7 = 8'hA8;
        i_im8 = 8'hB8;
        i_im9 = 8'hB6;
        #10 //3-20
        i_im1 = 8'h39;
        i_im2 = 8'h3B;
        i_im3 = 8'hB8;
        i_im4 = 8'h35;
        i_im5 = 8'hBB;
        i_im6 = 8'h20;
        i_im7 = 8'hB8;
        i_im8 = 8'hB6;
        i_im9 = 8'h33;
        #10 //3-21
        i_im1 = 8'h3B;
        i_im2 = 8'hB8;
        i_im3 = 8'h3B;
        i_im4 = 8'hBB;
        i_im5 = 8'h20;
        i_im6 = 8'h35;
        i_im7 = 8'hB6;
        i_im8 = 8'h33;
        i_im9 = 8'h3C;
        #10 //3-22
        i_im1 = 8'hB8;
        i_im2 = 8'h3B;
        i_im3 = 8'hAF;
        i_im4 = 8'h20;
        i_im5 = 8'h35;
        i_im6 = 8'hB9;
        i_im7 = 8'h33;
        i_im8 = 8'h3C;
        i_im9 = 8'hB9;
        #10 //3-23
        i_im1 = 8'h3B;
        i_im2 = 8'hAF;
        i_im3 = 8'hBA;
        i_im4 = 8'h35;
        i_im5 = 8'hB9;
        i_im6 = 8'h39;
        i_im7 = 8'h3C;
        i_im8 = 8'hB9;
        i_im9 = 8'h36;
        #10 //3-24
        i_im1 = 8'hAF;
        i_im2 = 8'hBA;
        i_im3 = 8'h38;
        i_im4 = 8'hB9;
        i_im5 = 8'h39;
        i_im6 = 8'hB1;
        i_im7 = 8'hB9;
        i_im8 = 8'h36;
        i_im9 = 8'hBA;
        #10 //3-25
        i_im1 = 8'hBA;
        i_im2 = 8'h38;
        i_im3 = 8'h2B;
        i_im4 = 8'h39;
        i_im5 = 8'hB1;
        i_im6 = 8'hBB;
        i_im7 = 8'h36;
        i_im8 = 8'hBA;
        i_im9 = 8'h38;
        #10 //3-26
        i_im1 = 8'h38;
        i_im2 = 8'h2B;
        i_im3 = 8'h34;
        i_im4 = 8'hB1;
        i_im5 = 8'hBB;
        i_im6 = 8'h30;
        i_im7 = 8'hBA;
        i_im8 = 8'h38;
        i_im9 = 8'hB6;
        #10 //4-1
        i_im1 = 8'hB4;
        i_im2 = 8'hB5;
        i_im3 = 8'hB9;
        i_im4 = 8'hBB;
        i_im5 = 8'h3A;
        i_im6 = 8'h39;
        i_im7 = 8'h39;
        i_im8 = 8'h3A;
        i_im9 = 8'hB5;
        #10 //4-2
        i_im1 = 8'hB5;
        i_im2 = 8'hB9;
        i_im3 = 8'hB7;
        i_im4 = 8'h3A;
        i_im5 = 8'h39;
        i_im6 = 8'h37;
        i_im7 = 8'h3A;
        i_im8 = 8'hB5;
        i_im9 = 8'h33;
        #10 //4-3
        i_im1 = 8'hB9;
        i_im2 = 8'hB7;
        i_im3 = 8'hB5;
        i_im4 = 8'h39;
        i_im5 = 8'h37;
        i_im6 = 8'hB7;
        i_im7 = 8'hB5;
        i_im8 = 8'h33;
        i_im9 = 8'hB2;
        #10 //4-4
        i_im1 = 8'hB7;
        i_im2 = 8'hB5;
        i_im3 = 8'hB7;
        i_im4 = 8'h37;
        i_im5 = 8'hB7;
        i_im6 = 8'h3A;
        i_im7 = 8'h33;
        i_im8 = 8'hB2;
        i_im9 = 8'hBA;
        #10 //4-5
        i_im1 = 8'hB5;
        i_im2 = 8'hB7;
        i_im3 = 8'hB4;
        i_im4 = 8'hB7;
        i_im5 = 8'h3A;
        i_im6 = 8'h20;
        i_im7 = 8'hB2;
        i_im8 = 8'hBA;
        i_im9 = 8'h3A;
        #10 //4-6
        i_im1 = 8'hB7;
        i_im2 = 8'hB4;
        i_im3 = 8'h3A;
        i_im4 = 8'h3A;
        i_im5 = 8'h20;
        i_im6 = 8'hBB;
        i_im7 = 8'hBA;
        i_im8 = 8'h3A;
        i_im9 = 8'hB8;
        #10 //4-7
        i_im1 = 8'hB4;
        i_im2 = 8'h3A;
        i_im3 = 8'hBB;
        i_im4 = 8'h20;
        i_im5 = 8'hBB;
        i_im6 = 8'hB9;
        i_im7 = 8'h3A;
        i_im8 = 8'hB8;
        i_im9 = 8'hBA;
        #10 //4-8
        i_im1 = 8'h3A;
        i_im2 = 8'hBB;
        i_im3 = 8'hB8;
        i_im4 = 8'hBB;
        i_im5 = 8'hB9;
        i_im6 = 8'h29;
        i_im7 = 8'hB8;
        i_im8 = 8'hBA;
        i_im9 = 8'hB4;
        #10 //4-9
        i_im1 = 8'hBB;
        i_im2 = 8'hB8;
        i_im3 = 8'hB1;
        i_im4 = 8'hB9;
        i_im5 = 8'h29;
        i_im6 = 8'hB8;
        i_im7 = 8'hBA;
        i_im8 = 8'hB4;
        i_im9 = 8'h36;
        #10 //4-10
        i_im1 = 8'hB8;
        i_im2 = 8'hB1;
        i_im3 = 8'hB2;
        i_im4 = 8'h29;
        i_im5 = 8'hB8;
        i_im6 = 8'hB1;
        i_im7 = 8'hB4;
        i_im8 = 8'h36;
        i_im9 = 8'h3A;
        #10 //4-11
        i_im1 = 8'hB1;
        i_im2 = 8'hB2;
        i_im3 = 8'hB2;
        i_im4 = 8'hB8;
        i_im5 = 8'hB1;
        i_im6 = 8'hA5;
        i_im7 = 8'h36;
        i_im8 = 8'h3A;
        i_im9 = 8'h30;
        #10 //4-12
        i_im1 = 8'hB2;
        i_im2 = 8'hB2;
        i_im3 = 8'hB8;
        i_im4 = 8'hB1;
        i_im5 = 8'hA5;
        i_im6 = 8'hBA;
        i_im7 = 8'h3A;
        i_im8 = 8'h30;
        i_im9 = 8'h3B;
        #10 //4-13
        i_im1 = 8'hB2;
        i_im2 = 8'hB8;
        i_im3 = 8'h39;
        i_im4 = 8'hA5;
        i_im5 = 8'hBA;
        i_im6 = 8'hBA;
        i_im7 = 8'h30;
        i_im8 = 8'h3B;
        i_im9 = 8'hBB;
        #10 //4-14
        i_im1 = 8'hB8;
        i_im2 = 8'h39;
        i_im3 = 8'h39;
        i_im4 = 8'hBA;
        i_im5 = 8'hBA;
        i_im6 = 8'h30;
        i_im7 = 8'h3B;
        i_im8 = 8'hBB;
        i_im9 = 8'hBA;
        #10 //4-15
        i_im1 = 8'h39;
        i_im2 = 8'h39;
        i_im3 = 8'hBB;
        i_im4 = 8'hBA;
        i_im5 = 8'h30;
        i_im6 = 8'h36;
        i_im7 = 8'hBB;
        i_im8 = 8'hBA;
        i_im9 = 8'h39;
        #10 //4-16
        i_im1 = 8'h39;
        i_im2 = 8'hBB;
        i_im3 = 8'hB7;
        i_im4 = 8'h30;
        i_im5 = 8'h36;
        i_im6 = 8'hB9;
        i_im7 = 8'hBA;
        i_im8 = 8'h39;
        i_im9 = 8'hAC;
        #10 //4-17
        i_im1 = 8'hBB;
        i_im2 = 8'hB7;
        i_im3 = 8'h35;
        i_im4 = 8'h36;
        i_im5 = 8'hB9;
        i_im6 = 8'hA8;
        i_im7 = 8'h39;
        i_im8 = 8'hAC;
        i_im9 = 8'hAD;
        #10 //4-18
        i_im1 = 8'hB7;
        i_im2 = 8'h35;
        i_im3 = 8'h35;
        i_im4 = 8'hB9;
        i_im5 = 8'hA8;
        i_im6 = 8'hB8;
        i_im7 = 8'hAC;
        i_im8 = 8'hAD;
        i_im9 = 8'hBB;
        #10 //4-19
        i_im1 = 8'h35;
        i_im2 = 8'h35;
        i_im3 = 8'hBB;
        i_im4 = 8'hA8;
        i_im5 = 8'hB8;
        i_im6 = 8'hB6;
        i_im7 = 8'hAD;
        i_im8 = 8'hBB;
        i_im9 = 8'hAE;
        #10 //4-20
        i_im1 = 8'h35;
        i_im2 = 8'hBB;
        i_im3 = 8'h20;
        i_im4 = 8'hB8;
        i_im5 = 8'hB6;
        i_im6 = 8'h33;
        i_im7 = 8'hBB;
        i_im8 = 8'hAE;
        i_im9 = 8'hB8;
        #10 //4-21
        i_im1 = 8'hBB;
        i_im2 = 8'h20;
        i_im3 = 8'h35;
        i_im4 = 8'hB6;
        i_im5 = 8'h33;
        i_im6 = 8'h3C;
        i_im7 = 8'hAE;
        i_im8 = 8'hB8;
        i_im9 = 8'hB0;
        #10 //4-22
        i_im1 = 8'h20;
        i_im2 = 8'h35;
        i_im3 = 8'hB9;
        i_im4 = 8'h33;
        i_im5 = 8'h3C;
        i_im6 = 8'hB9;
        i_im7 = 8'hB8;
        i_im8 = 8'hB0;
        i_im9 = 8'h37;
        #10 //4-23
        i_im1 = 8'h35;
        i_im2 = 8'hB9;
        i_im3 = 8'h39;
        i_im4 = 8'h3C;
        i_im5 = 8'hB9;
        i_im6 = 8'h36;
        i_im7 = 8'hB0;
        i_im8 = 8'h37;
        i_im9 = 8'h3B;
        #10 //4-24
        i_im1 = 8'hB9;
        i_im2 = 8'h39;
        i_im3 = 8'hB1;
        i_im4 = 8'hB9;
        i_im5 = 8'h36;
        i_im6 = 8'hBA;
        i_im7 = 8'h37;
        i_im8 = 8'h3B;
        i_im9 = 8'h37;
        #10 //4-25
        i_im1 = 8'h39;
        i_im2 = 8'hB1;
        i_im3 = 8'hBB;
        i_im4 = 8'h36;
        i_im5 = 8'hBA;
        i_im6 = 8'h38;
        i_im7 = 8'h3B;
        i_im8 = 8'h37;
        i_im9 = 8'h3B;
        #10 //4-26
        i_im1 = 8'hB1;
        i_im2 = 8'hBB;
        i_im3 = 8'h30;
        i_im4 = 8'hBA;
        i_im5 = 8'h38;
        i_im6 = 8'hB6;
        i_im7 = 8'h37;
        i_im8 = 8'h3B;
        i_im9 = 8'hBC;
        #10 //5-1
        i_im1 = 8'hBB;
        i_im2 = 8'h3A;
        i_im3 = 8'h39;
        i_im4 = 8'h39;
        i_im5 = 8'h3A;
        i_im6 = 8'hB5;
        i_im7 = 8'hBA;
        i_im8 = 8'hA7;
        i_im9 = 8'h35;
        #10 //5-2
        i_im1 = 8'h3A;
        i_im2 = 8'h39;
        i_im3 = 8'h37;
        i_im4 = 8'h3A;
        i_im5 = 8'hB5;
        i_im6 = 8'h33;
        i_im7 = 8'hA7;
        i_im8 = 8'h35;
        i_im9 = 8'hBA;
        #10 //5-3
        i_im1 = 8'h39;
        i_im2 = 8'h37;
        i_im3 = 8'hB7;
        i_im4 = 8'hB5;
        i_im5 = 8'h33;
        i_im6 = 8'hB2;
        i_im7 = 8'h35;
        i_im8 = 8'hBA;
        i_im9 = 8'h3A;
        #10 //5-4
        i_im1 = 8'h37;
        i_im2 = 8'hB7;
        i_im3 = 8'h3A;
        i_im4 = 8'h33;
        i_im5 = 8'hB2;
        i_im6 = 8'hBA;
        i_im7 = 8'hBA;
        i_im8 = 8'h3A;
        i_im9 = 8'h2E;
        #10 //5-5
        i_im1 = 8'hB7;
        i_im2 = 8'h3A;
        i_im3 = 8'h20;
        i_im4 = 8'hB2;
        i_im5 = 8'hBA;
        i_im6 = 8'h3A;
        i_im7 = 8'h3A;
        i_im8 = 8'h2E;
        i_im9 = 8'h3A;
        #10 //5-6
        i_im1 = 8'h3A;
        i_im2 = 8'h20;
        i_im3 = 8'hBB;
        i_im4 = 8'hBA;
        i_im5 = 8'h3A;
        i_im6 = 8'hB8;
        i_im7 = 8'h2E;
        i_im8 = 8'h3A;
        i_im9 = 8'hB8;
        #10 //5-7
        i_im1 = 8'h20;
        i_im2 = 8'hBB;
        i_im3 = 8'hB9;
        i_im4 = 8'h3A;
        i_im5 = 8'hB8;
        i_im6 = 8'hBA;
        i_im7 = 8'h3A;
        i_im8 = 8'hB8;
        i_im9 = 8'h39;
        #10 //5-8
        i_im1 = 8'hBB;
        i_im2 = 8'hB9;
        i_im3 = 8'h29;
        i_im4 = 8'hB8;
        i_im5 = 8'hBA;
        i_im6 = 8'hB4;
        i_im7 = 8'hB8;
        i_im8 = 8'h39;
        i_im9 = 8'h3B;
        #10 //5-9
        i_im1 = 8'hB9;
        i_im2 = 8'h29;
        i_im3 = 8'hB8;
        i_im4 = 8'hBA;
        i_im5 = 8'hB4;
        i_im6 = 8'h36;
        i_im7 = 8'h39;
        i_im8 = 8'h3B;
        i_im9 = 8'hB6;
        #10 //5-10
        i_im1 = 8'h29;
        i_im2 = 8'hB8;
        i_im3 = 8'hB1;
        i_im4 = 8'hB4;
        i_im5 = 8'h36;
        i_im6 = 8'h3A;
        i_im7 = 8'h3B;
        i_im8 = 8'hB6;
        i_im9 = 8'hB6;
        #10 //5-11
        i_im1 = 8'hB8;
        i_im2 = 8'hB1;
        i_im3 = 8'hA5;
        i_im4 = 8'h36;
        i_im5 = 8'h3A;
        i_im6 = 8'h30;
        i_im7 = 8'hB6;
        i_im8 = 8'hB6;
        i_im9 = 8'hB9;
        #10 //5-12
        i_im1 = 8'hB1;
        i_im2 = 8'hA5;
        i_im3 = 8'hBA;
        i_im4 = 8'h3A;
        i_im5 = 8'h30;
        i_im6 = 8'h3B;
        i_im7 = 8'hB6;
        i_im8 = 8'hB9;
        i_im9 = 8'h3A;
        #10 //5-13
        i_im1 = 8'hA5;
        i_im2 = 8'hBA;
        i_im3 = 8'hBA;
        i_im4 = 8'h30;
        i_im5 = 8'h3B;
        i_im6 = 8'hBB;
        i_im7 = 8'hB9;
        i_im8 = 8'h3A;
        i_im9 = 8'hAE;
        #10 //5-14
        i_im1 = 8'hBA;
        i_im2 = 8'hBA;
        i_im3 = 8'h30;
        i_im4 = 8'h3B;
        i_im5 = 8'hBB;
        i_im6 = 8'hBA;
        i_im7 = 8'h3A;
        i_im8 = 8'hAE;
        i_im9 = 8'h31;
        #10 //5-15
        i_im1 = 8'hBA;
        i_im2 = 8'h30;
        i_im3 = 8'h36;
        i_im4 = 8'hBB;
        i_im5 = 8'hBA;
        i_im6 = 8'h39;
        i_im7 = 8'hAE;
        i_im8 = 8'h31;
        i_im9 = 8'hB1;
        #10 //5-16
        i_im1 = 8'h30;
        i_im2 = 8'h36;
        i_im3 = 8'hB9;
        i_im4 = 8'hBA;
        i_im5 = 8'h39;
        i_im6 = 8'hAC;
        i_im7 = 8'h31;
        i_im8 = 8'hB1;
        i_im9 = 8'hB6;
        #10 //5-17
        i_im1 = 8'h36;
        i_im2 = 8'hB9;
        i_im3 = 8'hA8;
        i_im4 = 8'h39;
        i_im5 = 8'hAC;
        i_im6 = 8'hAD;
        i_im7 = 8'hB1;
        i_im8 = 8'hB6;
        i_im9 = 8'h39;
        #10 //5-18
        i_im1 = 8'hB9;
        i_im2 = 8'hA8;
        i_im3 = 8'hB8;
        i_im4 = 8'hAC;
        i_im5 = 8'hAD;
        i_im6 = 8'hBB;
        i_im7 = 8'hB6;
        i_im8 = 8'h39;
        i_im9 = 8'hB7;
        #10 //5-19
        i_im1 = 8'hA8;
        i_im2 = 8'hB8;
        i_im3 = 8'hB6;
        i_im4 = 8'hAD;
        i_im5 = 8'hBB;
        i_im6 = 8'hAE;
        i_im7 = 8'h39;
        i_im8 = 8'hB7;
        i_im9 = 8'hB6;
        #10 //5-20
        i_im1 = 8'hB8;
        i_im2 = 8'hB6;
        i_im3 = 8'h33;
        i_im4 = 8'hBB;
        i_im5 = 8'hAE;
        i_im6 = 8'hB8;
        i_im7 = 8'hB7;
        i_im8 = 8'hB6;
        i_im9 = 8'h35;
        #10 //5-21
        i_im1 = 8'hB6;
        i_im2 = 8'h33;
        i_im3 = 8'h3C;
        i_im4 = 8'hAE;
        i_im5 = 8'hB8;
        i_im6 = 8'hB0;
        i_im7 = 8'hB6;
        i_im8 = 8'h35;
        i_im9 = 8'hB9;
        #10 //5-22
        i_im1 = 8'h33;
        i_im2 = 8'h3C;
        i_im3 = 8'hB9;
        i_im4 = 8'hB8;
        i_im5 = 8'hB0;
        i_im6 = 8'h37;
        i_im7 = 8'h35;
        i_im8 = 8'hB9;
        i_im9 = 8'hB8;
        #10 //5-23
        i_im1 = 8'h3C;
        i_im2 = 8'hB9;
        i_im3 = 8'h36;
        i_im4 = 8'hB0;
        i_im5 = 8'h37;
        i_im6 = 8'h3B;
        i_im7 = 8'hB9;
        i_im8 = 8'hB8;
        i_im9 = 8'hB5;
        #10 //5-24
        i_im1 = 8'hB9;
        i_im2 = 8'h36;
        i_im3 = 8'hBA;
        i_im4 = 8'h37;
        i_im5 = 8'h3B;
        i_im6 = 8'h37;
        i_im7 = 8'hB8;
        i_im8 = 8'hB5;
        i_im9 = 8'hA6;
        #10 //5-25
        i_im1 = 8'h36;
        i_im2 = 8'hBA;
        i_im3 = 8'h38;
        i_im4 = 8'h3B;
        i_im5 = 8'h37;
        i_im6 = 8'h3B;
        i_im7 = 8'hB5;
        i_im8 = 8'hA6;
        i_im9 = 8'hB1;
        #10 //5-26
        i_im1 = 8'hBA;
        i_im2 = 8'h38;
        i_im3 = 8'hB6;
        i_im4 = 8'h37;
        i_im5 = 8'h3B;
        i_im6 = 8'hBC;
        i_im7 = 8'hA6;
        i_im8 = 8'hB1;
        i_im9 = 8'h39;
        #10 //6-1
        i_im1 = 8'h39;
        i_im2 = 8'h3A;
        i_im3 = 8'hB5;
        i_im4 = 8'hBA;
        i_im5 = 8'hA7;
        i_im6 = 8'h35;
        i_im7 = 8'h34;
        i_im8 = 8'hBA;
        i_im9 = 8'h35;
        #10 //6-2
        i_im1 = 8'h3A;
        i_im2 = 8'hB5;
        i_im3 = 8'h33;
        i_im4 = 8'hA7;
        i_im5 = 8'h35;
        i_im6 = 8'hBA;
        i_im7 = 8'hBA;
        i_im8 = 8'h35;
        i_im9 = 8'h3C;
        #10 //6-3
        i_im1 = 8'hB5;
        i_im2 = 8'h33;
        i_im3 = 8'hB2;
        i_im4 = 8'h35;
        i_im5 = 8'hBA;
        i_im6 = 8'h3A;
        i_im7 = 8'h35;
        i_im8 = 8'h3C;
        i_im9 = 8'h3B;
        #10 //6-4
        i_im1 = 8'h33;
        i_im2 = 8'hB2;
        i_im3 = 8'hBA;
        i_im4 = 8'hBA;
        i_im5 = 8'h3A;
        i_im6 = 8'h2E;
        i_im7 = 8'h3C;
        i_im8 = 8'h3B;
        i_im9 = 8'hB5;
        #10 //6-5
        i_im1 = 8'hB2;
        i_im2 = 8'hBA;
        i_im3 = 8'h3A;
        i_im4 = 8'h3A;
        i_im5 = 8'h2E;
        i_im6 = 8'h3A;
        i_im7 = 8'h3B;
        i_im8 = 8'hB5;
        i_im9 = 8'h38;
        #10 //6-6
        i_im1 = 8'hBA;
        i_im2 = 8'h3A;
        i_im3 = 8'hB8;
        i_im4 = 8'h2E;
        i_im5 = 8'h3A;
        i_im6 = 8'hB8;
        i_im7 = 8'hB5;
        i_im8 = 8'h38;
        i_im9 = 8'hBA;
        #10 //6-7
        i_im1 = 8'h3A;
        i_im2 = 8'hB8;
        i_im3 = 8'hBA;
        i_im4 = 8'h3A;
        i_im5 = 8'hB8;
        i_im6 = 8'h39;
        i_im7 = 8'h38;
        i_im8 = 8'hBA;
        i_im9 = 8'hB7;
        #10 //6-8
        i_im1 = 8'hB8;
        i_im2 = 8'hBA;
        i_im3 = 8'hB4;
        i_im4 = 8'hB8;
        i_im5 = 8'h39;
        i_im6 = 8'h3B;
        i_im7 = 8'hBA;
        i_im8 = 8'hB7;
        i_im9 = 8'h1C;
        #10 //6-9
        i_im1 = 8'hBA;
        i_im2 = 8'hB4;
        i_im3 = 8'h36;
        i_im4 = 8'h39;
        i_im5 = 8'h3B;
        i_im6 = 8'hB6;
        i_im7 = 8'hB7;
        i_im8 = 8'h1C;
        i_im9 = 8'h34;
        #10 //6-10
        i_im1 = 8'hB4;
        i_im2 = 8'h36;
        i_im3 = 8'h3A;
        i_im4 = 8'h3B;
        i_im5 = 8'hB6;
        i_im6 = 8'hB6;
        i_im7 = 8'h1C;
        i_im8 = 8'h34;
        i_im9 = 8'hB9;
        #10 //6-11
        i_im1 = 8'h36;
        i_im2 = 8'h3A;
        i_im3 = 8'h30;
        i_im4 = 8'hB6;
        i_im5 = 8'hB6;
        i_im6 = 8'hB9;
        i_im7 = 8'h34;
        i_im8 = 8'hB9;
        i_im9 = 8'h38;
        #10 //6-12
        i_im1 = 8'h3A;
        i_im2 = 8'h30;
        i_im3 = 8'h3B;
        i_im4 = 8'hB6;
        i_im5 = 8'hB9;
        i_im6 = 8'h3A;
        i_im7 = 8'hB9;
        i_im8 = 8'h38;
        i_im9 = 8'h2F;
        #10 //6-13
        i_im1 = 8'h30;
        i_im2 = 8'h3B;
        i_im3 = 8'hBB;
        i_im4 = 8'hB9;
        i_im5 = 8'h3A;
        i_im6 = 8'hAE;
        i_im7 = 8'h38;
        i_im8 = 8'h2F;
        i_im9 = 8'hAE;
        #10 //6-14
        i_im1 = 8'h3B;
        i_im2 = 8'hBB;
        i_im3 = 8'hBA;
        i_im4 = 8'h3A;
        i_im5 = 8'hAE;
        i_im6 = 8'h31;
        i_im7 = 8'h2F;
        i_im8 = 8'hAE;
        i_im9 = 8'h3A;
        #10 //6-15
        i_im1 = 8'hBB;
        i_im2 = 8'hBA;
        i_im3 = 8'h39;
        i_im4 = 8'hAE;
        i_im5 = 8'h31;
        i_im6 = 8'hB1;
        i_im7 = 8'hAE;
        i_im8 = 8'h3A;
        i_im9 = 8'h37;
        #10 //6-16
        i_im1 = 8'hBA;
        i_im2 = 8'h39;
        i_im3 = 8'hAC;
        i_im4 = 8'h31;
        i_im5 = 8'hB1;
        i_im6 = 8'hB6;
        i_im7 = 8'h3A;
        i_im8 = 8'h37;
        i_im9 = 8'hBB;
        #10 //6-17
        i_im1 = 8'h39;
        i_im2 = 8'hAC;
        i_im3 = 8'hAD;
        i_im4 = 8'hB1;
        i_im5 = 8'hB6;
        i_im6 = 8'h39;
        i_im7 = 8'h37;
        i_im8 = 8'hBB;
        i_im9 = 8'hB9;
        #10 //6-18
        i_im1 = 8'hAC;
        i_im2 = 8'hAD;
        i_im3 = 8'hBB;
        i_im4 = 8'hB6;
        i_im5 = 8'h39;
        i_im6 = 8'hB7;
        i_im7 = 8'hBB;
        i_im8 = 8'hB9;
        i_im9 = 8'h39;
        #10 //6-19
        i_im1 = 8'hAD;
        i_im2 = 8'hBB;
        i_im3 = 8'hAE;
        i_im4 = 8'h39;
        i_im5 = 8'hB7;
        i_im6 = 8'hB6;
        i_im7 = 8'hB9;
        i_im8 = 8'h39;
        i_im9 = 8'h39;
        #10 //6-20
        i_im1 = 8'hBB;
        i_im2 = 8'hAE;
        i_im3 = 8'hB8;
        i_im4 = 8'hB7;
        i_im5 = 8'hB6;
        i_im6 = 8'h35;
        i_im7 = 8'h39;
        i_im8 = 8'h39;
        i_im9 = 8'hB6;
        #10 //6-21
        i_im1 = 8'hAE;
        i_im2 = 8'hB8;
        i_im3 = 8'hB0;
        i_im4 = 8'hB6;
        i_im5 = 8'h35;
        i_im6 = 8'hB9;
        i_im7 = 8'h39;
        i_im8 = 8'hB6;
        i_im9 = 8'hB8;
        #10 //6-22
        i_im1 = 8'hB8;
        i_im2 = 8'hB0;
        i_im3 = 8'h37;
        i_im4 = 8'h35;
        i_im5 = 8'hB9;
        i_im6 = 8'hB8;
        i_im7 = 8'hB6;
        i_im8 = 8'hB8;
        i_im9 = 8'hA9;
        #10 //6-23
        i_im1 = 8'hB0;
        i_im2 = 8'h37;
        i_im3 = 8'h3B;
        i_im4 = 8'hB9;
        i_im5 = 8'hB8;
        i_im6 = 8'hB5;
        i_im7 = 8'hB8;
        i_im8 = 8'hA9;
        i_im9 = 8'h2C;
        #10 //6-24
        i_im1 = 8'h37;
        i_im2 = 8'h3B;
        i_im3 = 8'h37;
        i_im4 = 8'hB8;
        i_im5 = 8'hB5;
        i_im6 = 8'hA6;
        i_im7 = 8'hA9;
        i_im8 = 8'h2C;
        i_im9 = 8'h38;
        #10 //6-25
        i_im1 = 8'h3B;
        i_im2 = 8'h37;
        i_im3 = 8'h3B;
        i_im4 = 8'hB5;
        i_im5 = 8'hA6;
        i_im6 = 8'hB1;
        i_im7 = 8'h2C;
        i_im8 = 8'h38;
        i_im9 = 8'hBC;
        #10 //6-26
        i_im1 = 8'h37;
        i_im2 = 8'h3B;
        i_im3 = 8'hBC;
        i_im4 = 8'hA6;
        i_im5 = 8'hB1;
        i_im6 = 8'h39;
        i_im7 = 8'h38;
        i_im8 = 8'hBC;
        i_im9 = 8'h3B;
        #10 //7-1
        i_im1 = 8'hBA;
        i_im2 = 8'hA7;
        i_im3 = 8'h35;
        i_im4 = 8'h34;
        i_im5 = 8'hBA;
        i_im6 = 8'h35;
        i_im7 = 8'h34;
        i_im8 = 8'h2D;
        i_im9 = 8'hB6;
        #10 //7-2
        i_im1 = 8'hA7;
        i_im2 = 8'h35;
        i_im3 = 8'hBA;
        i_im4 = 8'hBA;
        i_im5 = 8'h35;
        i_im6 = 8'h3C;
        i_im7 = 8'h2D;
        i_im8 = 8'hB6;
        i_im9 = 8'hBC;
        #10 //7-3
        i_im1 = 8'h35;
        i_im2 = 8'hBA;
        i_im3 = 8'h3A;
        i_im4 = 8'h35;
        i_im5 = 8'h3C;
        i_im6 = 8'h3B;
        i_im7 = 8'hB6;
        i_im8 = 8'hBC;
        i_im9 = 8'hA7;
        #10 //7-4
        i_im1 = 8'hBA;
        i_im2 = 8'h3A;
        i_im3 = 8'h2E;
        i_im4 = 8'h3C;
        i_im5 = 8'h3B;
        i_im6 = 8'hB5;
        i_im7 = 8'hBC;
        i_im8 = 8'hA7;
        i_im9 = 8'hBA;
        #10 //7-5
        i_im1 = 8'h3A;
        i_im2 = 8'h2E;
        i_im3 = 8'h3A;
        i_im4 = 8'h3B;
        i_im5 = 8'hB5;
        i_im6 = 8'h38;
        i_im7 = 8'hA7;
        i_im8 = 8'hBA;
        i_im9 = 8'h35;
        #10 //7-6
        i_im1 = 8'h2E;
        i_im2 = 8'h3A;
        i_im3 = 8'hB8;
        i_im4 = 8'hB5;
        i_im5 = 8'h38;
        i_im6 = 8'hBA;
        i_im7 = 8'hBA;
        i_im8 = 8'h35;
        i_im9 = 8'hB4;
        #10 //7-7
        i_im1 = 8'h3A;
        i_im2 = 8'hB8;
        i_im3 = 8'h39;
        i_im4 = 8'h38;
        i_im5 = 8'hBA;
        i_im6 = 8'hB7;
        i_im7 = 8'h35;
        i_im8 = 8'hB4;
        i_im9 = 8'hB4;
        #10 //7-8
        i_im1 = 8'hB8;
        i_im2 = 8'h39;
        i_im3 = 8'h3B;
        i_im4 = 8'hBA;
        i_im5 = 8'hB7;
        i_im6 = 8'h1C;
        i_im7 = 8'hB4;
        i_im8 = 8'hB4;
        i_im9 = 8'hBA;
        #10 //7-9
        i_im1 = 8'h39;
        i_im2 = 8'h3B;
        i_im3 = 8'hB6;
        i_im4 = 8'hB7;
        i_im5 = 8'h1C;
        i_im6 = 8'h34;
        i_im7 = 8'hB4;
        i_im8 = 8'hBA;
        i_im9 = 8'hBC;
        #10 //7-10
        i_im1 = 8'h3B;
        i_im2 = 8'hB6;
        i_im3 = 8'hB6;
        i_im4 = 8'h1C;
        i_im5 = 8'h34;
        i_im6 = 8'hB9;
        i_im7 = 8'hBA;
        i_im8 = 8'hBC;
        i_im9 = 8'h34;
        #10 //7-11
        i_im1 = 8'hB6;
        i_im2 = 8'hB6;
        i_im3 = 8'hB9;
        i_im4 = 8'h34;
        i_im5 = 8'hB9;
        i_im6 = 8'h38;
        i_im7 = 8'hBC;
        i_im8 = 8'h34;
        i_im9 = 8'h3B;
        #10 //7-12
        i_im1 = 8'hB6;
        i_im2 = 8'hB9;
        i_im3 = 8'h3A;
        i_im4 = 8'hB9;
        i_im5 = 8'h38;
        i_im6 = 8'h2F;
        i_im7 = 8'h34;
        i_im8 = 8'h3B;
        i_im9 = 8'h2C;
        #10 //7-13
        i_im1 = 8'hB9;
        i_im2 = 8'h3A;
        i_im3 = 8'hAE;
        i_im4 = 8'h38;
        i_im5 = 8'h2F;
        i_im6 = 8'hAE;
        i_im7 = 8'h3B;
        i_im8 = 8'h2C;
        i_im9 = 8'hB7;
        #10 //7-14
        i_im1 = 8'h3A;
        i_im2 = 8'hAE;
        i_im3 = 8'h31;
        i_im4 = 8'h2F;
        i_im5 = 8'hAE;
        i_im6 = 8'h3A;
        i_im7 = 8'h2C;
        i_im8 = 8'hB7;
        i_im9 = 8'h2C;
        #10 //7-15
        i_im1 = 8'hAE;
        i_im2 = 8'h31;
        i_im3 = 8'hB1;
        i_im4 = 8'hAE;
        i_im5 = 8'h3A;
        i_im6 = 8'h37;
        i_im7 = 8'hB7;
        i_im8 = 8'h2C;
        i_im9 = 8'hBC;
        #10 //7-16
        i_im1 = 8'h31;
        i_im2 = 8'hB1;
        i_im3 = 8'hB6;
        i_im4 = 8'h3A;
        i_im5 = 8'h37;
        i_im6 = 8'hBB;
        i_im7 = 8'h2C;
        i_im8 = 8'hBC;
        i_im9 = 8'hB9;
        #10 //7-17
        i_im1 = 8'hB1;
        i_im2 = 8'hB6;
        i_im3 = 8'h39;
        i_im4 = 8'h37;
        i_im5 = 8'hBB;
        i_im6 = 8'hB9;
        i_im7 = 8'hBC;
        i_im8 = 8'hB9;
        i_im9 = 8'h3A;
        #10 //7-18
        i_im1 = 8'hB6;
        i_im2 = 8'h39;
        i_im3 = 8'hB7;
        i_im4 = 8'hBB;
        i_im5 = 8'hB9;
        i_im6 = 8'h39;
        i_im7 = 8'hB9;
        i_im8 = 8'h3A;
        i_im9 = 8'hBB;
        #10 //7-19
        i_im1 = 8'h39;
        i_im2 = 8'hB7;
        i_im3 = 8'hB6;
        i_im4 = 8'hB9;
        i_im5 = 8'h39;
        i_im6 = 8'h39;
        i_im7 = 8'h3A;
        i_im8 = 8'hBB;
        i_im9 = 8'h3B;
        #10 //7-20
        i_im1 = 8'hB7;
        i_im2 = 8'hB6;
        i_im3 = 8'h35;
        i_im4 = 8'h39;
        i_im5 = 8'h39;
        i_im6 = 8'hB6;
        i_im7 = 8'hBB;
        i_im8 = 8'h3B;
        i_im9 = 8'hB4;
        #10 //7-21
        i_im1 = 8'hB6;
        i_im2 = 8'h35;
        i_im3 = 8'hB9;
        i_im4 = 8'h39;
        i_im5 = 8'hB6;
        i_im6 = 8'hB8;
        i_im7 = 8'h3B;
        i_im8 = 8'hB4;
        i_im9 = 8'hB5;
        #10 //7-22
        i_im1 = 8'h35;
        i_im2 = 8'hB9;
        i_im3 = 8'hB8;
        i_im4 = 8'hB6;
        i_im5 = 8'hB8;
        i_im6 = 8'hA9;
        i_im7 = 8'hB4;
        i_im8 = 8'hB5;
        i_im9 = 8'h3A;
        #10 //7-23
        i_im1 = 8'hB9;
        i_im2 = 8'hB8;
        i_im3 = 8'hB5;
        i_im4 = 8'hB8;
        i_im5 = 8'hA9;
        i_im6 = 8'h2C;
        i_im7 = 8'hB5;
        i_im8 = 8'h3A;
        i_im9 = 8'h3B;
        #10 //7-24
        i_im1 = 8'hB8;
        i_im2 = 8'hB5;
        i_im3 = 8'hA6;
        i_im4 = 8'hA9;
        i_im5 = 8'h2C;
        i_im6 = 8'h38;
        i_im7 = 8'h3A;
        i_im8 = 8'h3B;
        i_im9 = 8'hAE;
        #10 //7-25
        i_im1 = 8'hB5;
        i_im2 = 8'hA6;
        i_im3 = 8'hB1;
        i_im4 = 8'h2C;
        i_im5 = 8'h38;
        i_im6 = 8'hBC;
        i_im7 = 8'h3B;
        i_im8 = 8'hAE;
        i_im9 = 8'hA5;
        #10 //7-26
        i_im1 = 8'hA6;
        i_im2 = 8'hB1;
        i_im3 = 8'h39;
        i_im4 = 8'h38;
        i_im5 = 8'hBC;
        i_im6 = 8'h3B;
        i_im7 = 8'hAE;
        i_im8 = 8'hA5;
        i_im9 = 8'h3B;
        #10 //8-1
        i_im1 = 8'h34;
        i_im2 = 8'hBA;
        i_im3 = 8'h35;
        i_im4 = 8'h34;
        i_im5 = 8'h2D;
        i_im6 = 8'hB6;
        i_im7 = 8'h33;
        i_im8 = 8'h35;
        i_im9 = 8'h32;
        #10 //8-2
        i_im1 = 8'hBA;
        i_im2 = 8'h35;
        i_im3 = 8'h3C;
        i_im4 = 8'h2D;
        i_im5 = 8'hB6;
        i_im6 = 8'hBC;
        i_im7 = 8'h35;
        i_im8 = 8'h32;
        i_im9 = 8'h39;
        #10 //8-3
        i_im1 = 8'h35;
        i_im2 = 8'h3C;
        i_im3 = 8'h3B;
        i_im4 = 8'hB6;
        i_im5 = 8'hBC;
        i_im6 = 8'hA7;
        i_im7 = 8'h32;
        i_im8 = 8'h39;
        i_im9 = 8'hB7;
        #10 //8-4
        i_im1 = 8'h3C;
        i_im2 = 8'h3B;
        i_im3 = 8'hB5;
        i_im4 = 8'hBC;
        i_im5 = 8'hA7;
        i_im6 = 8'hBA;
        i_im7 = 8'h39;
        i_im8 = 8'hB7;
        i_im9 = 8'hB8;
        #10 //8-5
        i_im1 = 8'h3B;
        i_im2 = 8'hB5;
        i_im3 = 8'h38;
        i_im4 = 8'hA7;
        i_im5 = 8'hBA;
        i_im6 = 8'h35;
        i_im7 = 8'hB7;
        i_im8 = 8'hB8;
        i_im9 = 8'h35;
        #10 //8-6
        i_im1 = 8'hB5;
        i_im2 = 8'h38;
        i_im3 = 8'hBA;
        i_im4 = 8'hBA;
        i_im5 = 8'h35;
        i_im6 = 8'hB4;
        i_im7 = 8'hB8;
        i_im8 = 8'h35;
        i_im9 = 8'h38;
        #10 //8-7
        i_im1 = 8'h38;
        i_im2 = 8'hBA;
        i_im3 = 8'hB7;
        i_im4 = 8'h35;
        i_im5 = 8'hB4;
        i_im6 = 8'hB4;
        i_im7 = 8'h35;
        i_im8 = 8'h38;
        i_im9 = 8'h36;
        #10 //8-8
        i_im1 = 8'hBA;
        i_im2 = 8'hB7;
        i_im3 = 8'h1C;
        i_im4 = 8'hB4;
        i_im5 = 8'hB4;
        i_im6 = 8'hBA;
        i_im7 = 8'h38;
        i_im8 = 8'h36;
        i_im9 = 8'h3C;
        #10 //8-9
        i_im1 = 8'hB7;
        i_im2 = 8'h1C;
        i_im3 = 8'h34;
        i_im4 = 8'hB4;
        i_im5 = 8'hBA;
        i_im6 = 8'hBC;
        i_im7 = 8'h36;
        i_im8 = 8'h3C;
        i_im9 = 8'hAC;
        #10 //8-10
        i_im1 = 8'h1C;
        i_im2 = 8'h34;
        i_im3 = 8'hB9;
        i_im4 = 8'hBA;
        i_im5 = 8'hBC;
        i_im6 = 8'h34;
        i_im7 = 8'h3C;
        i_im8 = 8'hAC;
        i_im9 = 8'h29;
        #10 //8-11
        i_im1 = 8'h34;
        i_im2 = 8'hB9;
        i_im3 = 8'h38;
        i_im4 = 8'hBC;
        i_im5 = 8'h34;
        i_im6 = 8'h3B;
        i_im7 = 8'hAC;
        i_im8 = 8'h29;
        i_im9 = 8'hB9;
        #10 //8-12
        i_im1 = 8'hB9;
        i_im2 = 8'h38;
        i_im3 = 8'h2F;
        i_im4 = 8'h34;
        i_im5 = 8'h3B;
        i_im6 = 8'h2C;
        i_im7 = 8'h29;
        i_im8 = 8'hB9;
        i_im9 = 8'h39;
        #10 //8-13
        i_im1 = 8'h38;
        i_im2 = 8'h2F;
        i_im3 = 8'hAE;
        i_im4 = 8'h3B;
        i_im5 = 8'h2C;
        i_im6 = 8'hB7;
        i_im7 = 8'hB9;
        i_im8 = 8'h39;
        i_im9 = 8'h36;
        #10 //8-14
        i_im1 = 8'h2F;
        i_im2 = 8'hAE;
        i_im3 = 8'h3A;
        i_im4 = 8'h2C;
        i_im5 = 8'hB7;
        i_im6 = 8'h2C;
        i_im7 = 8'h39;
        i_im8 = 8'h36;
        i_im9 = 8'hBC;
        #10 //8-15
        i_im1 = 8'hAE;
        i_im2 = 8'h3A;
        i_im3 = 8'h37;
        i_im4 = 8'hB7;
        i_im5 = 8'h2C;
        i_im6 = 8'hBC;
        i_im7 = 8'h36;
        i_im8 = 8'hBC;
        i_im9 = 8'h3C;
        #10 //8-16
        i_im1 = 8'h3A;
        i_im2 = 8'h37;
        i_im3 = 8'hBB;
        i_im4 = 8'h2C;
        i_im5 = 8'hBC;
        i_im6 = 8'hB9;
        i_im7 = 8'hBC;
        i_im8 = 8'h3C;
        i_im9 = 8'hB7;
        #10 //8-17
        i_im1 = 8'h37;
        i_im2 = 8'hBB;
        i_im3 = 8'hB9;
        i_im4 = 8'hBC;
        i_im5 = 8'hB9;
        i_im6 = 8'h3A;
        i_im7 = 8'h3C;
        i_im8 = 8'hB7;
        i_im9 = 8'hAF;
        #10 //8-18
        i_im1 = 8'hBB;
        i_im2 = 8'hB9;
        i_im3 = 8'h39;
        i_im4 = 8'hB9;
        i_im5 = 8'h3A;
        i_im6 = 8'hBB;
        i_im7 = 8'hB7;
        i_im8 = 8'hAF;
        i_im9 = 8'h20;
        #10 //8-19
        i_im1 = 8'hB9;
        i_im2 = 8'h39;
        i_im3 = 8'h39;
        i_im4 = 8'h3A;
        i_im5 = 8'hBB;
        i_im6 = 8'h3B;
        i_im7 = 8'hAF;
        i_im8 = 8'h20;
        i_im9 = 8'h35;
        #10 //8-20
        i_im1 = 8'h39;
        i_im2 = 8'h39;
        i_im3 = 8'hB6;
        i_im4 = 8'hBB;
        i_im5 = 8'h3B;
        i_im6 = 8'hB4;
        i_im7 = 8'h20;
        i_im8 = 8'h35;
        i_im9 = 8'hBC;
        #10 //8-21
        i_im1 = 8'h39;
        i_im2 = 8'hB6;
        i_im3 = 8'hB8;
        i_im4 = 8'h3B;
        i_im5 = 8'hB4;
        i_im6 = 8'hB5;
        i_im7 = 8'h35;
        i_im8 = 8'hBC;
        i_im9 = 8'hBB;
        #10 //8-22
        i_im1 = 8'hB6;
        i_im2 = 8'hB8;
        i_im3 = 8'hA9;
        i_im4 = 8'hB4;
        i_im5 = 8'hB5;
        i_im6 = 8'h3A;
        i_im7 = 8'hBC;
        i_im8 = 8'hBB;
        i_im9 = 8'h3B;
        #10 //8-23
        i_im1 = 8'hB8;
        i_im2 = 8'hA9;
        i_im3 = 8'h2C;
        i_im4 = 8'hB5;
        i_im5 = 8'h3A;
        i_im6 = 8'h3B;
        i_im7 = 8'hBB;
        i_im8 = 8'h3B;
        i_im9 = 8'hB7;
        #10 //8-24
        i_im1 = 8'hA9;
        i_im2 = 8'h2C;
        i_im3 = 8'h38;
        i_im4 = 8'h3A;
        i_im5 = 8'h3B;
        i_im6 = 8'hAE;
        i_im7 = 8'h3B;
        i_im8 = 8'hB7;
        i_im9 = 8'hAC;
        #10 //8-25
        i_im1 = 8'h2C;
        i_im2 = 8'h38;
        i_im3 = 8'hBC;
        i_im4 = 8'h3B;
        i_im5 = 8'hAE;
        i_im6 = 8'hA5;
        i_im7 = 8'hB7;
        i_im8 = 8'hAC;
        i_im9 = 8'h3B;
        #10 //8-26
        i_im1 = 8'h38;
        i_im2 = 8'hBC;
        i_im3 = 8'h3B;
        i_im4 = 8'hAE;
        i_im5 = 8'hA5;
        i_im6 = 8'h3B;
        i_im7 = 8'hAC;
        i_im8 = 8'h3B;
        i_im9 = 8'h2E;
        #10 //9-1
        i_im1 = 8'h34;
        i_im2 = 8'h2D;
        i_im3 = 8'hB6;
        i_im4 = 8'h33;
        i_im5 = 8'h35;
        i_im6 = 8'h32;
        i_im7 = 8'hB1;
        i_im8 = 8'h39;
        i_im9 = 8'hB5;
        #10 //9-2
        i_im1 = 8'h2D;
        i_im2 = 8'hB6;
        i_im3 = 8'hBC;
        i_im4 = 8'h35;
        i_im5 = 8'h32;
        i_im6 = 8'h39;
        i_im7 = 8'h39;
        i_im8 = 8'hB5;
        i_im9 = 8'h38;
        #10 //9-3
        i_im1 = 8'hB6;
        i_im2 = 8'hBC;
        i_im3 = 8'hA7;
        i_im4 = 8'h32;
        i_im5 = 8'h39;
        i_im6 = 8'hB7;
        i_im7 = 8'hB5;
        i_im8 = 8'h38;
        i_im9 = 8'h20;
        #10 //9-4
        i_im1 = 8'hBC;
        i_im2 = 8'hA7;
        i_im3 = 8'hBA;
        i_im4 = 8'h39;
        i_im5 = 8'hB7;
        i_im6 = 8'hB8;
        i_im7 = 8'h38;
        i_im8 = 8'h20;
        i_im9 = 8'h3B;
        #10 //9-5
        i_im1 = 8'hA7;
        i_im2 = 8'hBA;
        i_im3 = 8'h35;
        i_im4 = 8'hB7;
        i_im5 = 8'hB8;
        i_im6 = 8'h35;
        i_im7 = 8'h20;
        i_im8 = 8'h3B;
        i_im9 = 8'hBA;
        #10 //9-6
        i_im1 = 8'hBA;
        i_im2 = 8'h35;
        i_im3 = 8'hB4;
        i_im4 = 8'hB8;
        i_im5 = 8'h35;
        i_im6 = 8'h38;
        i_im7 = 8'h3B;
        i_im8 = 8'hBA;
        i_im9 = 8'h32;
        #10 //9-7
        i_im1 = 8'h35;
        i_im2 = 8'hB4;
        i_im3 = 8'hB4;
        i_im4 = 8'h35;
        i_im5 = 8'h38;
        i_im6 = 8'h36;
        i_im7 = 8'hBA;
        i_im8 = 8'h32;
        i_im9 = 8'h32;
        #10 //9-8
        i_im1 = 8'hB4;
        i_im2 = 8'hB4;
        i_im3 = 8'hBA;
        i_im4 = 8'h38;
        i_im5 = 8'h36;
        i_im6 = 8'h3C;
        i_im7 = 8'h32;
        i_im8 = 8'h32;
        i_im9 = 8'hBA;
        #10 //9-9
        i_im1 = 8'hB4;
        i_im2 = 8'hBA;
        i_im3 = 8'hBC;
        i_im4 = 8'h36;
        i_im5 = 8'h3C;
        i_im6 = 8'hAC;
        i_im7 = 8'h32;
        i_im8 = 8'hBA;
        i_im9 = 8'hAF;
        #10 //9-10
        i_im1 = 8'hBA;
        i_im2 = 8'hBC;
        i_im3 = 8'h34;
        i_im4 = 8'h3C;
        i_im5 = 8'hAC;
        i_im6 = 8'h29;
        i_im7 = 8'hBA;
        i_im8 = 8'hAF;
        i_im9 = 8'h39;
        #10 //9-11
        i_im1 = 8'hBC;
        i_im2 = 8'h34;
        i_im3 = 8'h3B;
        i_im4 = 8'hAC;
        i_im5 = 8'h29;
        i_im6 = 8'hB9;
        i_im7 = 8'hAF;
        i_im8 = 8'h39;
        i_im9 = 8'h39;
        #10 //9-12
        i_im1 = 8'h34;
        i_im2 = 8'h3B;
        i_im3 = 8'h2C;
        i_im4 = 8'h29;
        i_im5 = 8'hB9;
        i_im6 = 8'h39;
        i_im7 = 8'h39;
        i_im8 = 8'h39;
        i_im9 = 8'h26;
        #10 //9-13
        i_im1 = 8'h3B;
        i_im2 = 8'h2C;
        i_im3 = 8'hB7;
        i_im4 = 8'hB9;
        i_im5 = 8'h39;
        i_im6 = 8'h36;
        i_im7 = 8'h39;
        i_im8 = 8'h26;
        i_im9 = 8'h39;
        #10 //9-14
        i_im1 = 8'h2C;
        i_im2 = 8'hB7;
        i_im3 = 8'h2C;
        i_im4 = 8'h39;
        i_im5 = 8'h36;
        i_im6 = 8'hBC;
        i_im7 = 8'h26;
        i_im8 = 8'h39;
        i_im9 = 8'hB6;
        #10 //9-15
        i_im1 = 8'hB7;
        i_im2 = 8'h2C;
        i_im3 = 8'hBC;
        i_im4 = 8'h36;
        i_im5 = 8'hBC;
        i_im6 = 8'h3C;
        i_im7 = 8'h39;
        i_im8 = 8'hB6;
        i_im9 = 8'h3C;
        #10 //9-16
        i_im1 = 8'h2C;
        i_im2 = 8'hBC;
        i_im3 = 8'hB9;
        i_im4 = 8'hBC;
        i_im5 = 8'h3C;
        i_im6 = 8'hB7;
        i_im7 = 8'hB6;
        i_im8 = 8'h3C;
        i_im9 = 8'h2A;
        #10 //9-17
        i_im1 = 8'hBC;
        i_im2 = 8'hB9;
        i_im3 = 8'h3A;
        i_im4 = 8'h3C;
        i_im5 = 8'hB7;
        i_im6 = 8'hAF;
        i_im7 = 8'h3C;
        i_im8 = 8'h2A;
        i_im9 = 8'hB7;
        #10 //9-18
        i_im1 = 8'hB9;
        i_im2 = 8'h3A;
        i_im3 = 8'hBB;
        i_im4 = 8'hB7;
        i_im5 = 8'hAF;
        i_im6 = 8'h20;
        i_im7 = 8'h2A;
        i_im8 = 8'hB7;
        i_im9 = 8'h39;
        #10 //9-19
        i_im1 = 8'h3A;
        i_im2 = 8'hBB;
        i_im3 = 8'h3B;
        i_im4 = 8'hAF;
        i_im5 = 8'h20;
        i_im6 = 8'h35;
        i_im7 = 8'hB7;
        i_im8 = 8'h39;
        i_im9 = 8'h37;
        #10 //9-20
        i_im1 = 8'hBB;
        i_im2 = 8'h3B;
        i_im3 = 8'hB4;
        i_im4 = 8'h20;
        i_im5 = 8'h35;
        i_im6 = 8'hBC;
        i_im7 = 8'h39;
        i_im8 = 8'h37;
        i_im9 = 8'h36;
        #10 //9-21
        i_im1 = 8'h3B;
        i_im2 = 8'hB4;
        i_im3 = 8'hB5;
        i_im4 = 8'h35;
        i_im5 = 8'hBC;
        i_im6 = 8'hBB;
        i_im7 = 8'h37;
        i_im8 = 8'h36;
        i_im9 = 8'h38;
        #10 //9-22
        i_im1 = 8'hB4;
        i_im2 = 8'hB5;
        i_im3 = 8'h3A;
        i_im4 = 8'hBC;
        i_im5 = 8'hBB;
        i_im6 = 8'h3B;
        i_im7 = 8'h36;
        i_im8 = 8'h38;
        i_im9 = 8'h36;
        #10 //9-23
        i_im1 = 8'hB5;
        i_im2 = 8'h3A;
        i_im3 = 8'h3B;
        i_im4 = 8'hBB;
        i_im5 = 8'h3B;
        i_im6 = 8'hB7;
        i_im7 = 8'h38;
        i_im8 = 8'h36;
        i_im9 = 8'hBC;
        #10 //9-24
        i_im1 = 8'h3A;
        i_im2 = 8'h3B;
        i_im3 = 8'hAE;
        i_im4 = 8'h3B;
        i_im5 = 8'hB7;
        i_im6 = 8'hAC;
        i_im7 = 8'h36;
        i_im8 = 8'hBC;
        i_im9 = 8'h37;
        #10 //9-25
        i_im1 = 8'h3B;
        i_im2 = 8'hAE;
        i_im3 = 8'hA5;
        i_im4 = 8'hB7;
        i_im5 = 8'hAC;
        i_im6 = 8'h3B;
        i_im7 = 8'hBC;
        i_im8 = 8'h37;
        i_im9 = 8'hBB;
        #10 //9-26
        i_im1 = 8'hAE;
        i_im2 = 8'hA5;
        i_im3 = 8'h3B;
        i_im4 = 8'hAC;
        i_im5 = 8'h3B;
        i_im6 = 8'h2E;
        i_im7 = 8'h37;
        i_im8 = 8'hBB;
        i_im9 = 8'h36;
        #10 //10-1
        i_im1 = 8'h33;
        i_im2 = 8'h35;
        i_im3 = 8'h32;
        i_im4 = 8'hB1;
        i_im5 = 8'h39;
        i_im6 = 8'hB5;
        i_im7 = 8'h39;
        i_im8 = 8'h3B;
        i_im9 = 8'hB9;
        #10 //10-2
        i_im1 = 8'h35;
        i_im2 = 8'h32;
        i_im3 = 8'h39;
        i_im4 = 8'h39;
        i_im5 = 8'hB5;
        i_im6 = 8'h38;
        i_im7 = 8'h3B;
        i_im8 = 8'hB9;
        i_im9 = 8'hBA;
        #10 //10-3
        i_im1 = 8'h32;
        i_im2 = 8'h39;
        i_im3 = 8'hB7;
        i_im4 = 8'hB5;
        i_im5 = 8'h38;
        i_im6 = 8'h20;
        i_im7 = 8'hB9;
        i_im8 = 8'hBA;
        i_im9 = 8'hB9;
        #10 //10-4
        i_im1 = 8'h39;
        i_im2 = 8'hB7;
        i_im3 = 8'hB8;
        i_im4 = 8'h38;
        i_im5 = 8'h20;
        i_im6 = 8'h3B;
        i_im7 = 8'hBA;
        i_im8 = 8'hB9;
        i_im9 = 8'hB5;
        #10 //10-5
        i_im1 = 8'hB7;
        i_im2 = 8'hB8;
        i_im3 = 8'h35;
        i_im4 = 8'h20;
        i_im5 = 8'h3B;
        i_im6 = 8'hBA;
        i_im7 = 8'hB9;
        i_im8 = 8'hB5;
        i_im9 = 8'hBB;
        #10 //10-6
        i_im1 = 8'hB8;
        i_im2 = 8'h35;
        i_im3 = 8'h38;
        i_im4 = 8'h3B;
        i_im5 = 8'hBA;
        i_im6 = 8'h32;
        i_im7 = 8'hB5;
        i_im8 = 8'hBB;
        i_im9 = 8'hB4;
        #10 //10-7
        i_im1 = 8'h35;
        i_im2 = 8'h38;
        i_im3 = 8'h36;
        i_im4 = 8'hBA;
        i_im5 = 8'h32;
        i_im6 = 8'h32;
        i_im7 = 8'hBB;
        i_im8 = 8'hB4;
        i_im9 = 8'h38;
        #10 //10-8
        i_im1 = 8'h38;
        i_im2 = 8'h36;
        i_im3 = 8'h3C;
        i_im4 = 8'h32;
        i_im5 = 8'h32;
        i_im6 = 8'hBA;
        i_im7 = 8'hB4;
        i_im8 = 8'h38;
        i_im9 = 8'hBC;
        #10 //10-9
        i_im1 = 8'h36;
        i_im2 = 8'h3C;
        i_im3 = 8'hAC;
        i_im4 = 8'h32;
        i_im5 = 8'hBA;
        i_im6 = 8'hAF;
        i_im7 = 8'h38;
        i_im8 = 8'hBC;
        i_im9 = 8'hB9;
        #10 //10-10
        i_im1 = 8'h3C;
        i_im2 = 8'hAC;
        i_im3 = 8'h29;
        i_im4 = 8'hBA;
        i_im5 = 8'hAF;
        i_im6 = 8'h39;
        i_im7 = 8'hBC;
        i_im8 = 8'hB9;
        i_im9 = 8'h33;
        #10 //10-11
        i_im1 = 8'hAC;
        i_im2 = 8'h29;
        i_im3 = 8'hB9;
        i_im4 = 8'hAF;
        i_im5 = 8'h39;
        i_im6 = 8'h39;
        i_im7 = 8'hB9;
        i_im8 = 8'h33;
        i_im9 = 8'hBB;
        #10 //10-12
        i_im1 = 8'h29;
        i_im2 = 8'hB9;
        i_im3 = 8'h39;
        i_im4 = 8'h39;
        i_im5 = 8'h39;
        i_im6 = 8'h26;
        i_im7 = 8'h33;
        i_im8 = 8'hBB;
        i_im9 = 8'hBC;
        #10 //10-13
        i_im1 = 8'hB9;
        i_im2 = 8'h39;
        i_im3 = 8'h36;
        i_im4 = 8'h39;
        i_im5 = 8'h26;
        i_im6 = 8'h39;
        i_im7 = 8'hBB;
        i_im8 = 8'hBC;
        i_im9 = 8'h30;
        #10 //10-14
        i_im1 = 8'h39;
        i_im2 = 8'h36;
        i_im3 = 8'hBC;
        i_im4 = 8'h26;
        i_im5 = 8'h39;
        i_im6 = 8'hB6;
        i_im7 = 8'hBC;
        i_im8 = 8'h30;
        i_im9 = 8'h36;
        #10 //10-15
        i_im1 = 8'h36;
        i_im2 = 8'hBC;
        i_im3 = 8'h3C;
        i_im4 = 8'h39;
        i_im5 = 8'hB6;
        i_im6 = 8'h3C;
        i_im7 = 8'h30;
        i_im8 = 8'h36;
        i_im9 = 8'h36;
        #10 //10-16
        i_im1 = 8'hBC;
        i_im2 = 8'h3C;
        i_im3 = 8'hB7;
        i_im4 = 8'hB6;
        i_im5 = 8'h3C;
        i_im6 = 8'h2A;
        i_im7 = 8'h36;
        i_im8 = 8'h36;
        i_im9 = 8'h3A;
        #10 //10-17
        i_im1 = 8'h3C;
        i_im2 = 8'hB7;
        i_im3 = 8'hAF;
        i_im4 = 8'h3C;
        i_im5 = 8'h2A;
        i_im6 = 8'hB7;
        i_im7 = 8'h36;
        i_im8 = 8'h3A;
        i_im9 = 8'hB8;
        #10 //10-18
        i_im1 = 8'hB7;
        i_im2 = 8'hAF;
        i_im3 = 8'h20;
        i_im4 = 8'h2A;
        i_im5 = 8'hB7;
        i_im6 = 8'h39;
        i_im7 = 8'h3A;
        i_im8 = 8'hB8;
        i_im9 = 8'hB8;
        #10 //10-19
        i_im1 = 8'hAF;
        i_im2 = 8'h20;
        i_im3 = 8'h35;
        i_im4 = 8'hB7;
        i_im5 = 8'h39;
        i_im6 = 8'h37;
        i_im7 = 8'hB8;
        i_im8 = 8'hB8;
        i_im9 = 8'h35;
        #10 //10-20
        i_im1 = 8'h20;
        i_im2 = 8'h35;
        i_im3 = 8'hBC;
        i_im4 = 8'h39;
        i_im5 = 8'h37;
        i_im6 = 8'h36;
        i_im7 = 8'hB8;
        i_im8 = 8'h35;
        i_im9 = 8'h36;
        #10 //10-21
        i_im1 = 8'h35;
        i_im2 = 8'hBC;
        i_im3 = 8'hBB;
        i_im4 = 8'h37;
        i_im5 = 8'h36;
        i_im6 = 8'h38;
        i_im7 = 8'h35;
        i_im8 = 8'h36;
        i_im9 = 8'hBC;
        #10 //10-22
        i_im1 = 8'hBC;
        i_im2 = 8'hBB;
        i_im3 = 8'h3B;
        i_im4 = 8'h36;
        i_im5 = 8'h38;
        i_im6 = 8'h36;
        i_im7 = 8'h36;
        i_im8 = 8'hBC;
        i_im9 = 8'h3C;
        #10 //10-23
        i_im1 = 8'hBB;
        i_im2 = 8'h3B;
        i_im3 = 8'hB7;
        i_im4 = 8'h38;
        i_im5 = 8'h36;
        i_im6 = 8'hBC;
        i_im7 = 8'hBC;
        i_im8 = 8'h3C;
        i_im9 = 8'h39;
        #10 //10-24
        i_im1 = 8'h3B;
        i_im2 = 8'hB7;
        i_im3 = 8'hAC;
        i_im4 = 8'h36;
        i_im5 = 8'hBC;
        i_im6 = 8'h37;
        i_im7 = 8'h3C;
        i_im8 = 8'h39;
        i_im9 = 8'h3B;
        #10 //10-25
        i_im1 = 8'hB7;
        i_im2 = 8'hAC;
        i_im3 = 8'h3B;
        i_im4 = 8'hBC;
        i_im5 = 8'h37;
        i_im6 = 8'hBB;
        i_im7 = 8'h39;
        i_im8 = 8'h3B;
        i_im9 = 8'h37;
        #10 //10-26
        i_im1 = 8'hAC;
        i_im2 = 8'h3B;
        i_im3 = 8'h2E;
        i_im4 = 8'h37;
        i_im5 = 8'hBB;
        i_im6 = 8'h36;
        i_im7 = 8'h3B;
        i_im8 = 8'h37;
        i_im9 = 8'h2B;
        #10 //11-1
        i_im1 = 8'hB1;
        i_im2 = 8'h39;
        i_im3 = 8'hB5;
        i_im4 = 8'h39;
        i_im5 = 8'h3B;
        i_im6 = 8'hB9;
        i_im7 = 8'hB7;
        i_im8 = 8'hB1;
        i_im9 = 8'hB5;
        #10 //11-2
        i_im1 = 8'h39;
        i_im2 = 8'hB5;
        i_im3 = 8'h38;
        i_im4 = 8'h3B;
        i_im5 = 8'hB9;
        i_im6 = 8'hBA;
        i_im7 = 8'hB1;
        i_im8 = 8'hB5;
        i_im9 = 8'h33;
        #10 //11-3
        i_im1 = 8'hB5;
        i_im2 = 8'h38;
        i_im3 = 8'h20;
        i_im4 = 8'hB9;
        i_im5 = 8'hBA;
        i_im6 = 8'hB9;
        i_im7 = 8'hB5;
        i_im8 = 8'h33;
        i_im9 = 8'h39;
        #10 //11-4
        i_im1 = 8'h38;
        i_im2 = 8'h20;
        i_im3 = 8'h3B;
        i_im4 = 8'hBA;
        i_im5 = 8'hB9;
        i_im6 = 8'hB5;
        i_im7 = 8'h33;
        i_im8 = 8'h39;
        i_im9 = 8'h39;
        #10 //11-5
        i_im1 = 8'h20;
        i_im2 = 8'h3B;
        i_im3 = 8'hBA;
        i_im4 = 8'hB9;
        i_im5 = 8'hB5;
        i_im6 = 8'hBB;
        i_im7 = 8'h39;
        i_im8 = 8'h39;
        i_im9 = 8'h29;
        #10 //11-6
        i_im1 = 8'h3B;
        i_im2 = 8'hBA;
        i_im3 = 8'h32;
        i_im4 = 8'hB5;
        i_im5 = 8'hBB;
        i_im6 = 8'hB4;
        i_im7 = 8'h39;
        i_im8 = 8'h29;
        i_im9 = 8'hBC;
        #10 //11-7
        i_im1 = 8'hBA;
        i_im2 = 8'h32;
        i_im3 = 8'h32;
        i_im4 = 8'hBB;
        i_im5 = 8'hB4;
        i_im6 = 8'h38;
        i_im7 = 8'h29;
        i_im8 = 8'hBC;
        i_im9 = 8'hBA;
        #10 //11-8
        i_im1 = 8'h32;
        i_im2 = 8'h32;
        i_im3 = 8'hBA;
        i_im4 = 8'hB4;
        i_im5 = 8'h38;
        i_im6 = 8'hBC;
        i_im7 = 8'hBC;
        i_im8 = 8'hBA;
        i_im9 = 8'h3A;
        #10 //11-9
        i_im1 = 8'h32;
        i_im2 = 8'hBA;
        i_im3 = 8'hAF;
        i_im4 = 8'h38;
        i_im5 = 8'hBC;
        i_im6 = 8'hB9;
        i_im7 = 8'hBA;
        i_im8 = 8'h3A;
        i_im9 = 8'hB2;
        #10 //11-10
        i_im1 = 8'hBA;
        i_im2 = 8'hAF;
        i_im3 = 8'h39;
        i_im4 = 8'hBC;
        i_im5 = 8'hB9;
        i_im6 = 8'h33;
        i_im7 = 8'h3A;
        i_im8 = 8'hB2;
        i_im9 = 8'hBA;
        #10 //11-11
        i_im1 = 8'hAF;
        i_im2 = 8'h39;
        i_im3 = 8'h39;
        i_im4 = 8'hB9;
        i_im5 = 8'h33;
        i_im6 = 8'hBB;
        i_im7 = 8'hB2;
        i_im8 = 8'hBA;
        i_im9 = 8'hAD;
        #10 //11-12
        i_im1 = 8'h39;
        i_im2 = 8'h39;
        i_im3 = 8'h26;
        i_im4 = 8'h33;
        i_im5 = 8'hBB;
        i_im6 = 8'hBC;
        i_im7 = 8'hBA;
        i_im8 = 8'hAD;
        i_im9 = 8'hB4;
        #10 //11-13
        i_im1 = 8'h39;
        i_im2 = 8'h26;
        i_im3 = 8'h39;
        i_im4 = 8'hBB;
        i_im5 = 8'hBC;
        i_im6 = 8'h30;
        i_im7 = 8'hAD;
        i_im8 = 8'hB4;
        i_im9 = 8'hB9;
        #10 //11-14
        i_im1 = 8'h26;
        i_im2 = 8'h39;
        i_im3 = 8'hB6;
        i_im4 = 8'hBC;
        i_im5 = 8'h30;
        i_im6 = 8'h36;
        i_im7 = 8'hB4;
        i_im8 = 8'hB9;
        i_im9 = 8'hB5;
        #10 //11-15
        i_im1 = 8'h39;
        i_im2 = 8'hB6;
        i_im3 = 8'h3C;
        i_im4 = 8'h30;
        i_im5 = 8'h36;
        i_im6 = 8'h36;
        i_im7 = 8'hB9;
        i_im8 = 8'hB5;
        i_im9 = 8'hB6;
        #10 //11-16
        i_im1 = 8'hB6;
        i_im2 = 8'h3C;
        i_im3 = 8'h2A;
        i_im4 = 8'h36;
        i_im5 = 8'h36;
        i_im6 = 8'h3A;
        i_im7 = 8'hB5;
        i_im8 = 8'hB6;
        i_im9 = 8'h33;
        #10 //11-17
        i_im1 = 8'h3C;
        i_im2 = 8'h2A;
        i_im3 = 8'hB7;
        i_im4 = 8'h36;
        i_im5 = 8'h3A;
        i_im6 = 8'hB8;
        i_im7 = 8'hB6;
        i_im8 = 8'h33;
        i_im9 = 8'hB9;
        #10 //11-18
        i_im1 = 8'h2A;
        i_im2 = 8'hB7;
        i_im3 = 8'h39;
        i_im4 = 8'h3A;
        i_im5 = 8'hB8;
        i_im6 = 8'hB8;
        i_im7 = 8'h33;
        i_im8 = 8'hB9;
        i_im9 = 8'h36;
        #10 //11-19
        i_im1 = 8'hB7;
        i_im2 = 8'h39;
        i_im3 = 8'h37;
        i_im4 = 8'hB8;
        i_im5 = 8'hB8;
        i_im6 = 8'h35;
        i_im7 = 8'hB9;
        i_im8 = 8'h36;
        i_im9 = 8'h3A;
        #10 //11-20
        i_im1 = 8'h39;
        i_im2 = 8'h37;
        i_im3 = 8'h36;
        i_im4 = 8'hB8;
        i_im5 = 8'h35;
        i_im6 = 8'h36;
        i_im7 = 8'h36;
        i_im8 = 8'h3A;
        i_im9 = 8'hBB;
        #10 //11-21
        i_im1 = 8'h37;
        i_im2 = 8'h36;
        i_im3 = 8'h38;
        i_im4 = 8'h35;
        i_im5 = 8'h36;
        i_im6 = 8'hBC;
        i_im7 = 8'h3A;
        i_im8 = 8'hBB;
        i_im9 = 8'hAC;
        #10 //11-22
        i_im1 = 8'h36;
        i_im2 = 8'h38;
        i_im3 = 8'h36;
        i_im4 = 8'h36;
        i_im5 = 8'hBC;
        i_im6 = 8'h3C;
        i_im7 = 8'hBB;
        i_im8 = 8'hAC;
        i_im9 = 8'hBA;
        #10 //11-23
        i_im1 = 8'h38;
        i_im2 = 8'h36;
        i_im3 = 8'hBC;
        i_im4 = 8'hBC;
        i_im5 = 8'h3C;
        i_im6 = 8'h39;
        i_im7 = 8'hAC;
        i_im8 = 8'hBA;
        i_im9 = 8'hB7;
        #10 //11-24
        i_im1 = 8'h36;
        i_im2 = 8'hBC;
        i_im3 = 8'h37;
        i_im4 = 8'h3C;
        i_im5 = 8'h39;
        i_im6 = 8'h3B;
        i_im7 = 8'hBA;
        i_im8 = 8'hB7;
        i_im9 = 8'h34;
        #10 //11-25
        i_im1 = 8'hBC;
        i_im2 = 8'h37;
        i_im3 = 8'hBB;
        i_im4 = 8'h39;
        i_im5 = 8'h3B;
        i_im6 = 8'h37;
        i_im7 = 8'hB7;
        i_im8 = 8'h34;
        i_im9 = 8'hBA;
        #10 //11-26
        i_im1 = 8'h37;
        i_im2 = 8'hBB;
        i_im3 = 8'h36;
        i_im4 = 8'h3B;
        i_im5 = 8'h37;
        i_im6 = 8'h2B;
        i_im7 = 8'h34;
        i_im8 = 8'hBA;
        i_im9 = 8'hBB;
        #10 //12-1
        i_im1 = 8'h39;
        i_im2 = 8'h3B;
        i_im3 = 8'hB9;
        i_im4 = 8'hB7;
        i_im5 = 8'hB1;
        i_im6 = 8'hB5;
        i_im7 = 8'h3A;
        i_im8 = 8'hB8;
        i_im9 = 8'h3C;
        #10 //12-2
        i_im1 = 8'h3B;
        i_im2 = 8'hB9;
        i_im3 = 8'hBA;
        i_im4 = 8'hB1;
        i_im5 = 8'hB5;
        i_im6 = 8'h33;
        i_im7 = 8'hB8;
        i_im8 = 8'h3C;
        i_im9 = 8'hB9;
        #10 //12-3
        i_im1 = 8'hB9;
        i_im2 = 8'hBA;
        i_im3 = 8'hB9;
        i_im4 = 8'hB5;
        i_im5 = 8'h33;
        i_im6 = 8'h39;
        i_im7 = 8'h3C;
        i_im8 = 8'hB9;
        i_im9 = 8'hB4;
        #10 //12-4
        i_im1 = 8'hBA;
        i_im2 = 8'hB9;
        i_im3 = 8'hB5;
        i_im4 = 8'h33;
        i_im5 = 8'h39;
        i_im6 = 8'h39;
        i_im7 = 8'hB9;
        i_im8 = 8'hB4;
        i_im9 = 8'hB5;
        #10 //12-5
        i_im1 = 8'hB9;
        i_im2 = 8'hB5;
        i_im3 = 8'hBB;
        i_im4 = 8'h39;
        i_im5 = 8'h39;
        i_im6 = 8'h29;
        i_im7 = 8'hB4;
        i_im8 = 8'hB5;
        i_im9 = 8'hAE;
        #10 //12-6
        i_im1 = 8'hB5;
        i_im2 = 8'hBB;
        i_im3 = 8'hB4;
        i_im4 = 8'h39;
        i_im5 = 8'h29;
        i_im6 = 8'hBC;
        i_im7 = 8'hB5;
        i_im8 = 8'hAE;
        i_im9 = 8'h38;
        #10 //12-7
        i_im1 = 8'hBB;
        i_im2 = 8'hB4;
        i_im3 = 8'h38;
        i_im4 = 8'h29;
        i_im5 = 8'hBC;
        i_im6 = 8'hBA;
        i_im7 = 8'hAE;
        i_im8 = 8'h38;
        i_im9 = 8'hBB;
        #10 //12-8
        i_im1 = 8'hB4;
        i_im2 = 8'h38;
        i_im3 = 8'hBC;
        i_im4 = 8'hBC;
        i_im5 = 8'hBA;
        i_im6 = 8'h3A;
        i_im7 = 8'h38;
        i_im8 = 8'hBB;
        i_im9 = 8'h3C;
        #10 //12-9
        i_im1 = 8'h38;
        i_im2 = 8'hBC;
        i_im3 = 8'hB9;
        i_im4 = 8'hBA;
        i_im5 = 8'h3A;
        i_im6 = 8'hB2;
        i_im7 = 8'hBB;
        i_im8 = 8'h3C;
        i_im9 = 8'h39;
        #10 //12-10
        i_im1 = 8'hBC;
        i_im2 = 8'hB9;
        i_im3 = 8'h33;
        i_im4 = 8'h3A;
        i_im5 = 8'hB2;
        i_im6 = 8'hBA;
        i_im7 = 8'h3C;
        i_im8 = 8'h39;
        i_im9 = 8'hBB;
        #10 //12-11
        i_im1 = 8'hB9;
        i_im2 = 8'h33;
        i_im3 = 8'hBB;
        i_im4 = 8'hB2;
        i_im5 = 8'hBA;
        i_im6 = 8'hAD;
        i_im7 = 8'h39;
        i_im8 = 8'hBB;
        i_im9 = 8'hB6;
        #10 //12-12
        i_im1 = 8'h33;
        i_im2 = 8'hBB;
        i_im3 = 8'hBC;
        i_im4 = 8'hBA;
        i_im5 = 8'hAD;
        i_im6 = 8'hB4;
        i_im7 = 8'hBB;
        i_im8 = 8'hB6;
        i_im9 = 8'hB7;
        #10 //12-13
        i_im1 = 8'hBB;
        i_im2 = 8'hBC;
        i_im3 = 8'h30;
        i_im4 = 8'hAD;
        i_im5 = 8'hB4;
        i_im6 = 8'hB9;
        i_im7 = 8'hB6;
        i_im8 = 8'hB7;
        i_im9 = 8'h34;
        #10 //12-14
        i_im1 = 8'hBC;
        i_im2 = 8'h30;
        i_im3 = 8'h36;
        i_im4 = 8'hB4;
        i_im5 = 8'hB9;
        i_im6 = 8'hB5;
        i_im7 = 8'hB7;
        i_im8 = 8'h34;
        i_im9 = 8'hA4;
        #10 //12-15
        i_im1 = 8'h30;
        i_im2 = 8'h36;
        i_im3 = 8'h36;
        i_im4 = 8'hB9;
        i_im5 = 8'hB5;
        i_im6 = 8'hB6;
        i_im7 = 8'h34;
        i_im8 = 8'hA4;
        i_im9 = 8'hBB;
        #10 //12-16
        i_im1 = 8'h36;
        i_im2 = 8'h36;
        i_im3 = 8'h3A;
        i_im4 = 8'hB5;
        i_im5 = 8'hB6;
        i_im6 = 8'h33;
        i_im7 = 8'hA4;
        i_im8 = 8'hBB;
        i_im9 = 8'hB1;
        #10 //12-17
        i_im1 = 8'h36;
        i_im2 = 8'h3A;
        i_im3 = 8'hB8;
        i_im4 = 8'hB6;
        i_im5 = 8'h33;
        i_im6 = 8'hB9;
        i_im7 = 8'hBB;
        i_im8 = 8'hB1;
        i_im9 = 8'h37;
        #10 //12-18
        i_im1 = 8'h3A;
        i_im2 = 8'hB8;
        i_im3 = 8'hB8;
        i_im4 = 8'h33;
        i_im5 = 8'hB9;
        i_im6 = 8'h36;
        i_im7 = 8'hB1;
        i_im8 = 8'h37;
        i_im9 = 8'h3A;
        #10 //12-19
        i_im1 = 8'hB8;
        i_im2 = 8'hB8;
        i_im3 = 8'h35;
        i_im4 = 8'hB9;
        i_im5 = 8'h36;
        i_im6 = 8'h3A;
        i_im7 = 8'h37;
        i_im8 = 8'h3A;
        i_im9 = 8'h1C;
        #10 //12-20
        i_im1 = 8'hB8;
        i_im2 = 8'h35;
        i_im3 = 8'h36;
        i_im4 = 8'h36;
        i_im5 = 8'h3A;
        i_im6 = 8'hBB;
        i_im7 = 8'h3A;
        i_im8 = 8'h1C;
        i_im9 = 8'hBA;
        #10 //12-21
        i_im1 = 8'h35;
        i_im2 = 8'h36;
        i_im3 = 8'hBC;
        i_im4 = 8'h3A;
        i_im5 = 8'hBB;
        i_im6 = 8'hAC;
        i_im7 = 8'h1C;
        i_im8 = 8'hBA;
        i_im9 = 8'h3B;
        #10 //12-22
        i_im1 = 8'h36;
        i_im2 = 8'hBC;
        i_im3 = 8'h3C;
        i_im4 = 8'hBB;
        i_im5 = 8'hAC;
        i_im6 = 8'hBA;
        i_im7 = 8'hBA;
        i_im8 = 8'h3B;
        i_im9 = 8'h39;
        #10 //12-23
        i_im1 = 8'hBC;
        i_im2 = 8'h3C;
        i_im3 = 8'h39;
        i_im4 = 8'hAC;
        i_im5 = 8'hBA;
        i_im6 = 8'hB7;
        i_im7 = 8'h3B;
        i_im8 = 8'h39;
        i_im9 = 8'h30;
        #10 //12-24
        i_im1 = 8'h3C;
        i_im2 = 8'h39;
        i_im3 = 8'h3B;
        i_im4 = 8'hBA;
        i_im5 = 8'hB7;
        i_im6 = 8'h34;
        i_im7 = 8'h39;
        i_im8 = 8'h30;
        i_im9 = 8'hB6;
        #10 //12-25
        i_im1 = 8'h39;
        i_im2 = 8'h3B;
        i_im3 = 8'h37;
        i_im4 = 8'hB7;
        i_im5 = 8'h34;
        i_im6 = 8'hBA;
        i_im7 = 8'h30;
        i_im8 = 8'hB6;
        i_im9 = 8'h3C;
        #10 //12-26
        i_im1 = 8'h3B;
        i_im2 = 8'h37;
        i_im3 = 8'h2B;
        i_im4 = 8'h34;
        i_im5 = 8'hBA;
        i_im6 = 8'hBB;
        i_im7 = 8'hB6;
        i_im8 = 8'h3C;
        i_im9 = 8'hB7;
        #10 //13-1
        i_im1 = 8'hB7;
        i_im2 = 8'hB1;
        i_im3 = 8'hB5;
        i_im4 = 8'h3A;
        i_im5 = 8'hB8;
        i_im6 = 8'h3C;
        i_im7 = 8'hAC;
        i_im8 = 8'hB9;
        i_im9 = 8'h3A;
        #10 //13-2
        i_im1 = 8'hB1;
        i_im2 = 8'hB5;
        i_im3 = 8'h33;
        i_im4 = 8'hB8;
        i_im5 = 8'h3C;
        i_im6 = 8'hB9;
        i_im7 = 8'hB9;
        i_im8 = 8'h3A;
        i_im9 = 8'hB1;
        #10 //13-3
        i_im1 = 8'hB5;
        i_im2 = 8'h33;
        i_im3 = 8'h39;
        i_im4 = 8'h3C;
        i_im5 = 8'hB9;
        i_im6 = 8'hB4;
        i_im7 = 8'h3A;
        i_im8 = 8'hB1;
        i_im9 = 8'h34;
        #10 //13-4
        i_im1 = 8'h33;
        i_im2 = 8'h39;
        i_im3 = 8'h39;
        i_im4 = 8'hB9;
        i_im5 = 8'hB4;
        i_im6 = 8'hB5;
        i_im7 = 8'hB1;
        i_im8 = 8'h34;
        i_im9 = 8'h39;
        #10 //13-5
        i_im1 = 8'h39;
        i_im2 = 8'h39;
        i_im3 = 8'h29;
        i_im4 = 8'hB4;
        i_im5 = 8'hB5;
        i_im6 = 8'hAE;
        i_im7 = 8'h34;
        i_im8 = 8'h39;
        i_im9 = 8'hB6;
        #10 //13-6
        i_im1 = 8'h39;
        i_im2 = 8'h29;
        i_im3 = 8'hBC;
        i_im4 = 8'hB5;
        i_im5 = 8'hAE;
        i_im6 = 8'h38;
        i_im7 = 8'h39;
        i_im8 = 8'hB6;
        i_im9 = 8'h30;
        #10 //13-7
        i_im1 = 8'h29;
        i_im2 = 8'hBC;
        i_im3 = 8'hBA;
        i_im4 = 8'hAE;
        i_im5 = 8'h38;
        i_im6 = 8'hBB;
        i_im7 = 8'hB6;
        i_im8 = 8'h30;
        i_im9 = 8'hB4;
        #10 //13-8
        i_im1 = 8'hBC;
        i_im2 = 8'hBA;
        i_im3 = 8'h3A;
        i_im4 = 8'h38;
        i_im5 = 8'hBB;
        i_im6 = 8'h3C;
        i_im7 = 8'h30;
        i_im8 = 8'hB4;
        i_im9 = 8'h38;
        #10 //13-9
        i_im1 = 8'hBA;
        i_im2 = 8'h3A;
        i_im3 = 8'hB2;
        i_im4 = 8'hBB;
        i_im5 = 8'h3C;
        i_im6 = 8'h39;
        i_im7 = 8'hB4;
        i_im8 = 8'h38;
        i_im9 = 8'h34;
        #10 //13-10
        i_im1 = 8'h3A;
        i_im2 = 8'hB2;
        i_im3 = 8'hBA;
        i_im4 = 8'h3C;
        i_im5 = 8'h39;
        i_im6 = 8'hBB;
        i_im7 = 8'h38;
        i_im8 = 8'h34;
        i_im9 = 8'h3C;
        #10 //13-11
        i_im1 = 8'hB2;
        i_im2 = 8'hBA;
        i_im3 = 8'hAD;
        i_im4 = 8'h39;
        i_im5 = 8'hBB;
        i_im6 = 8'hB6;
        i_im7 = 8'h34;
        i_im8 = 8'h3C;
        i_im9 = 8'hBA;
        #10 //13-12
        i_im1 = 8'hBA;
        i_im2 = 8'hAD;
        i_im3 = 8'hB4;
        i_im4 = 8'hBB;
        i_im5 = 8'hB6;
        i_im6 = 8'hB7;
        i_im7 = 8'h3C;
        i_im8 = 8'hBA;
        i_im9 = 8'h34;
        #10 //13-13
        i_im1 = 8'hAD;
        i_im2 = 8'hB4;
        i_im3 = 8'hB9;
        i_im4 = 8'hB6;
        i_im5 = 8'hB7;
        i_im6 = 8'h34;
        i_im7 = 8'hBA;
        i_im8 = 8'h34;
        i_im9 = 8'h3A;
        #10 //13-14
        i_im1 = 8'hB4;
        i_im2 = 8'hB9;
        i_im3 = 8'hB5;
        i_im4 = 8'hB7;
        i_im5 = 8'h34;
        i_im6 = 8'hA4;
        i_im7 = 8'h34;
        i_im8 = 8'h3A;
        i_im9 = 8'h38;
        #10 //13-15
        i_im1 = 8'hB9;
        i_im2 = 8'hB5;
        i_im3 = 8'hB6;
        i_im4 = 8'h34;
        i_im5 = 8'hA4;
        i_im6 = 8'hBB;
        i_im7 = 8'h3A;
        i_im8 = 8'h38;
        i_im9 = 8'hB8;
        #10 //13-16
        i_im1 = 8'hB5;
        i_im2 = 8'hB6;
        i_im3 = 8'h33;
        i_im4 = 8'hA4;
        i_im5 = 8'hBB;
        i_im6 = 8'hB1;
        i_im7 = 8'h38;
        i_im8 = 8'hB8;
        i_im9 = 8'hB1;
        #10 //13-17
        i_im1 = 8'hB6;
        i_im2 = 8'h33;
        i_im3 = 8'hB9;
        i_im4 = 8'hBB;
        i_im5 = 8'hB1;
        i_im6 = 8'h37;
        i_im7 = 8'hB8;
        i_im8 = 8'hB1;
        i_im9 = 8'hB4;
        #10 //13-18
        i_im1 = 8'h33;
        i_im2 = 8'hB9;
        i_im3 = 8'h36;
        i_im4 = 8'hB1;
        i_im5 = 8'h37;
        i_im6 = 8'h3A;
        i_im7 = 8'hB1;
        i_im8 = 8'hB4;
        i_im9 = 8'h32;
        #10 //13-19
        i_im1 = 8'hB9;
        i_im2 = 8'h36;
        i_im3 = 8'h3A;
        i_im4 = 8'h37;
        i_im5 = 8'h3A;
        i_im6 = 8'h1C;
        i_im7 = 8'hB4;
        i_im8 = 8'h32;
        i_im9 = 8'h37;
        #10 //13-20
        i_im1 = 8'h36;
        i_im2 = 8'h3A;
        i_im3 = 8'hBB;
        i_im4 = 8'h3A;
        i_im5 = 8'h1C;
        i_im6 = 8'hBA;
        i_im7 = 8'h32;
        i_im8 = 8'h37;
        i_im9 = 8'h3A;
        #10 //13-21
        i_im1 = 8'h3A;
        i_im2 = 8'hBB;
        i_im3 = 8'hAC;
        i_im4 = 8'h1C;
        i_im5 = 8'hBA;
        i_im6 = 8'h3B;
        i_im7 = 8'h37;
        i_im8 = 8'h3A;
        i_im9 = 8'h2F;
        #10 //13-22
        i_im1 = 8'hBB;
        i_im2 = 8'hAC;
        i_im3 = 8'hBA;
        i_im4 = 8'hBA;
        i_im5 = 8'h3B;
        i_im6 = 8'h39;
        i_im7 = 8'h3A;
        i_im8 = 8'h2F;
        i_im9 = 8'h3B;
        #10 //13-23
        i_im1 = 8'hAC;
        i_im2 = 8'hBA;
        i_im3 = 8'hB7;
        i_im4 = 8'h3B;
        i_im5 = 8'h39;
        i_im6 = 8'h30;
        i_im7 = 8'h2F;
        i_im8 = 8'h3B;
        i_im9 = 8'h36;
        #10 //13-24
        i_im1 = 8'hBA;
        i_im2 = 8'hB7;
        i_im3 = 8'h34;
        i_im4 = 8'h39;
        i_im5 = 8'h30;
        i_im6 = 8'hB6;
        i_im7 = 8'h3B;
        i_im8 = 8'h36;
        i_im9 = 8'hBA;
        #10 //13-25
        i_im1 = 8'hB7;
        i_im2 = 8'h34;
        i_im3 = 8'hBA;
        i_im4 = 8'h30;
        i_im5 = 8'hB6;
        i_im6 = 8'h3C;
        i_im7 = 8'h36;
        i_im8 = 8'hBA;
        i_im9 = 8'h3A;
        #10 //13-26
        i_im1 = 8'h34;
        i_im2 = 8'hBA;
        i_im3 = 8'hBB;
        i_im4 = 8'hB6;
        i_im5 = 8'h3C;
        i_im6 = 8'hB7;
        i_im7 = 8'hBA;
        i_im8 = 8'h3A;
        i_im9 = 8'h34;
        #10 //14-1
        i_im1 = 8'h3A;
        i_im2 = 8'hB8;
        i_im3 = 8'h3C;
        i_im4 = 8'hAC;
        i_im5 = 8'hB9;
        i_im6 = 8'h3A;
        i_im7 = 8'h2B;
        i_im8 = 8'h3C;
        i_im9 = 8'h2F;
        #10 //14-2
        i_im1 = 8'hB8;
        i_im2 = 8'h3C;
        i_im3 = 8'hB9;
        i_im4 = 8'hB9;
        i_im5 = 8'h3A;
        i_im6 = 8'hB1;
        i_im7 = 8'h3C;
        i_im8 = 8'h2F;
        i_im9 = 8'h3A;
        #10 //14-3
        i_im1 = 8'h3C;
        i_im2 = 8'hB9;
        i_im3 = 8'hB4;
        i_im4 = 8'h3A;
        i_im5 = 8'hB1;
        i_im6 = 8'h34;
        i_im7 = 8'h2F;
        i_im8 = 8'h3A;
        i_im9 = 8'hB5;
        #10 //14-4
        i_im1 = 8'hB9;
        i_im2 = 8'hB4;
        i_im3 = 8'hB5;
        i_im4 = 8'hB1;
        i_im5 = 8'h34;
        i_im6 = 8'h39;
        i_im7 = 8'h3A;
        i_im8 = 8'hB5;
        i_im9 = 8'h31;
        #10 //14-5
        i_im1 = 8'hB4;
        i_im2 = 8'hB5;
        i_im3 = 8'hAE;
        i_im4 = 8'h34;
        i_im5 = 8'h39;
        i_im6 = 8'hB6;
        i_im7 = 8'hB5;
        i_im8 = 8'h31;
        i_im9 = 8'hB9;
        #10 //14-6
        i_im1 = 8'hB5;
        i_im2 = 8'hAE;
        i_im3 = 8'h38;
        i_im4 = 8'h39;
        i_im5 = 8'hB6;
        i_im6 = 8'h30;
        i_im7 = 8'h31;
        i_im8 = 8'hB9;
        i_im9 = 8'h2B;
        #10 //14-7
        i_im1 = 8'hAE;
        i_im2 = 8'h38;
        i_im3 = 8'hBB;
        i_im4 = 8'hB6;
        i_im5 = 8'h30;
        i_im6 = 8'hB4;
        i_im7 = 8'hB9;
        i_im8 = 8'h2B;
        i_im9 = 8'hB2;
        #10 //14-8
        i_im1 = 8'h38;
        i_im2 = 8'hBB;
        i_im3 = 8'h3C;
        i_im4 = 8'h30;
        i_im5 = 8'hB4;
        i_im6 = 8'h38;
        i_im7 = 8'h2B;
        i_im8 = 8'hB2;
        i_im9 = 8'hB9;
        #10 //14-9
        i_im1 = 8'hBB;
        i_im2 = 8'h3C;
        i_im3 = 8'h39;
        i_im4 = 8'hB4;
        i_im5 = 8'h38;
        i_im6 = 8'h34;
        i_im7 = 8'hB2;
        i_im8 = 8'hB9;
        i_im9 = 8'hB5;
        #10 //14-10
        i_im1 = 8'h3C;
        i_im2 = 8'h39;
        i_im3 = 8'hBB;
        i_im4 = 8'h38;
        i_im5 = 8'h34;
        i_im6 = 8'h3C;
        i_im7 = 8'hB9;
        i_im8 = 8'hB5;
        i_im9 = 8'hB8;
        #10 //14-11
        i_im1 = 8'h39;
        i_im2 = 8'hBB;
        i_im3 = 8'hB6;
        i_im4 = 8'h34;
        i_im5 = 8'h3C;
        i_im6 = 8'hBA;
        i_im7 = 8'hB5;
        i_im8 = 8'hB8;
        i_im9 = 8'hBA;
        #10 //14-12
        i_im1 = 8'hBB;
        i_im2 = 8'hB6;
        i_im3 = 8'hB7;
        i_im4 = 8'h3C;
        i_im5 = 8'hBA;
        i_im6 = 8'h34;
        i_im7 = 8'hB8;
        i_im8 = 8'hBA;
        i_im9 = 8'h32;
        #10 //14-13
        i_im1 = 8'hB6;
        i_im2 = 8'hB7;
        i_im3 = 8'h34;
        i_im4 = 8'hBA;
        i_im5 = 8'h34;
        i_im6 = 8'h3A;
        i_im7 = 8'hBA;
        i_im8 = 8'h32;
        i_im9 = 8'hB9;
        #10 //14-14
        i_im1 = 8'hB7;
        i_im2 = 8'h34;
        i_im3 = 8'hA4;
        i_im4 = 8'h34;
        i_im5 = 8'h3A;
        i_im6 = 8'h38;
        i_im7 = 8'h32;
        i_im8 = 8'hB9;
        i_im9 = 8'hBC;
        #10 //14-15
        i_im1 = 8'h34;
        i_im2 = 8'hA4;
        i_im3 = 8'hBB;
        i_im4 = 8'h3A;
        i_im5 = 8'h38;
        i_im6 = 8'hB8;
        i_im7 = 8'hB9;
        i_im8 = 8'hBC;
        i_im9 = 8'hB9;
        #10 //14-16
        i_im1 = 8'hA4;
        i_im2 = 8'hBB;
        i_im3 = 8'hB1;
        i_im4 = 8'h38;
        i_im5 = 8'hB8;
        i_im6 = 8'hB1;
        i_im7 = 8'hBC;
        i_im8 = 8'hB9;
        i_im9 = 8'hBC;
        #10 //14-17
        i_im1 = 8'hBB;
        i_im2 = 8'hB1;
        i_im3 = 8'h37;
        i_im4 = 8'hB8;
        i_im5 = 8'hB1;
        i_im6 = 8'hB4;
        i_im7 = 8'hB9;
        i_im8 = 8'hBC;
        i_im9 = 8'hB4;
        #10 //14-18
        i_im1 = 8'hB1;
        i_im2 = 8'h37;
        i_im3 = 8'h3A;
        i_im4 = 8'hB1;
        i_im5 = 8'hB4;
        i_im6 = 8'h32;
        i_im7 = 8'hBC;
        i_im8 = 8'hB4;
        i_im9 = 8'hA7;
        #10 //14-19
        i_im1 = 8'h37;
        i_im2 = 8'h3A;
        i_im3 = 8'h1C;
        i_im4 = 8'hB4;
        i_im5 = 8'h32;
        i_im6 = 8'h37;
        i_im7 = 8'hB4;
        i_im8 = 8'hA7;
        i_im9 = 8'h20;
        #10 //14-20
        i_im1 = 8'h3A;
        i_im2 = 8'h1C;
        i_im3 = 8'hBA;
        i_im4 = 8'h32;
        i_im5 = 8'h37;
        i_im6 = 8'h3A;
        i_im7 = 8'hA7;
        i_im8 = 8'h20;
        i_im9 = 8'h28;
        #10 //14-21
        i_im1 = 8'h1C;
        i_im2 = 8'hBA;
        i_im3 = 8'h3B;
        i_im4 = 8'h37;
        i_im5 = 8'h3A;
        i_im6 = 8'h2F;
        i_im7 = 8'h20;
        i_im8 = 8'h28;
        i_im9 = 8'hBA;
        #10 //14-22
        i_im1 = 8'hBA;
        i_im2 = 8'h3B;
        i_im3 = 8'h39;
        i_im4 = 8'h3A;
        i_im5 = 8'h2F;
        i_im6 = 8'h3B;
        i_im7 = 8'h28;
        i_im8 = 8'hBA;
        i_im9 = 8'hBA;
        #10 //14-23
        i_im1 = 8'h3B;
        i_im2 = 8'h39;
        i_im3 = 8'h30;
        i_im4 = 8'h2F;
        i_im5 = 8'h3B;
        i_im6 = 8'h36;
        i_im7 = 8'hBA;
        i_im8 = 8'hBA;
        i_im9 = 8'h3A;
        #10 //14-24
        i_im1 = 8'h39;
        i_im2 = 8'h30;
        i_im3 = 8'hB6;
        i_im4 = 8'h3B;
        i_im5 = 8'h36;
        i_im6 = 8'hBA;
        i_im7 = 8'hBA;
        i_im8 = 8'h3A;
        i_im9 = 8'h3B;
        #10 //14-25
        i_im1 = 8'h30;
        i_im2 = 8'hB6;
        i_im3 = 8'h3C;
        i_im4 = 8'h36;
        i_im5 = 8'hBA;
        i_im6 = 8'h3A;
        i_im7 = 8'h3A;
        i_im8 = 8'h3B;
        i_im9 = 8'h39;
        #10 //14-26
        i_im1 = 8'hB6;
        i_im2 = 8'h3C;
        i_im3 = 8'hB7;
        i_im4 = 8'hBA;
        i_im5 = 8'h3A;
        i_im6 = 8'h34;
        i_im7 = 8'h3B;
        i_im8 = 8'h39;
        i_im9 = 8'hB9;
        #10 //15-1
        i_im1 = 8'hAC;
        i_im2 = 8'hB9;
        i_im3 = 8'h3A;
        i_im4 = 8'h2B;
        i_im5 = 8'h3C;
        i_im6 = 8'h2F;
        i_im7 = 8'h39;
        i_im8 = 8'h36;
        i_im9 = 8'hB3;
        #10 //15-2
        i_im1 = 8'hB9;
        i_im2 = 8'h3A;
        i_im3 = 8'hB1;
        i_im4 = 8'h3C;
        i_im5 = 8'h2F;
        i_im6 = 8'h3A;
        i_im7 = 8'h36;
        i_im8 = 8'hB3;
        i_im9 = 8'hB3;
        #10 //15-3
        i_im1 = 8'h3A;
        i_im2 = 8'hB1;
        i_im3 = 8'h34;
        i_im4 = 8'h2F;
        i_im5 = 8'h3A;
        i_im6 = 8'hB5;
        i_im7 = 8'hB3;
        i_im8 = 8'hB3;
        i_im9 = 8'hBA;
        #10 //15-4
        i_im1 = 8'hB1;
        i_im2 = 8'h34;
        i_im3 = 8'h39;
        i_im4 = 8'h3A;
        i_im5 = 8'hB5;
        i_im6 = 8'h31;
        i_im7 = 8'hB3;
        i_im8 = 8'hBA;
        i_im9 = 8'hB9;
        #10 //15-5
        i_im1 = 8'h34;
        i_im2 = 8'h39;
        i_im3 = 8'hB6;
        i_im4 = 8'hB5;
        i_im5 = 8'h31;
        i_im6 = 8'hB9;
        i_im7 = 8'hBA;
        i_im8 = 8'hB9;
        i_im9 = 8'hB5;
        #10 //15-6
        i_im1 = 8'h39;
        i_im2 = 8'hB6;
        i_im3 = 8'h30;
        i_im4 = 8'h31;
        i_im5 = 8'hB9;
        i_im6 = 8'h2B;
        i_im7 = 8'hB9;
        i_im8 = 8'hB5;
        i_im9 = 8'h3A;
        #10 //15-7
        i_im1 = 8'hB6;
        i_im2 = 8'h30;
        i_im3 = 8'hB4;
        i_im4 = 8'hB9;
        i_im5 = 8'h2B;
        i_im6 = 8'hB2;
        i_im7 = 8'hB5;
        i_im8 = 8'h3A;
        i_im9 = 8'h2E;
        #10 //15-8
        i_im1 = 8'h30;
        i_im2 = 8'hB4;
        i_im3 = 8'h38;
        i_im4 = 8'h2B;
        i_im5 = 8'hB2;
        i_im6 = 8'hB9;
        i_im7 = 8'h3A;
        i_im8 = 8'h2E;
        i_im9 = 8'hB9;
        #10 //15-9
        i_im1 = 8'hB4;
        i_im2 = 8'h38;
        i_im3 = 8'h34;
        i_im4 = 8'hB2;
        i_im5 = 8'hB9;
        i_im6 = 8'hB5;
        i_im7 = 8'h2E;
        i_im8 = 8'hB9;
        i_im9 = 8'hBA;
        #10 //15-10
        i_im1 = 8'h38;
        i_im2 = 8'h34;
        i_im3 = 8'h3C;
        i_im4 = 8'hB9;
        i_im5 = 8'hB5;
        i_im6 = 8'hB8;
        i_im7 = 8'hB9;
        i_im8 = 8'hBA;
        i_im9 = 8'hB8;
        #10 //15-11
        i_im1 = 8'h34;
        i_im2 = 8'h3C;
        i_im3 = 8'hBA;
        i_im4 = 8'hB5;
        i_im5 = 8'hB8;
        i_im6 = 8'hBA;
        i_im7 = 8'hBA;
        i_im8 = 8'hB8;
        i_im9 = 8'h35;
        #10 //15-12
        i_im1 = 8'h3C;
        i_im2 = 8'hBA;
        i_im3 = 8'h34;
        i_im4 = 8'hB8;
        i_im5 = 8'hBA;
        i_im6 = 8'h32;
        i_im7 = 8'hB8;
        i_im8 = 8'h35;
        i_im9 = 8'h3A;
        #10 //15-13
        i_im1 = 8'hBA;
        i_im2 = 8'h34;
        i_im3 = 8'h3A;
        i_im4 = 8'hBA;
        i_im5 = 8'h32;
        i_im6 = 8'hB9;
        i_im7 = 8'h35;
        i_im8 = 8'h3A;
        i_im9 = 8'h39;
        #10 //15-14
        i_im1 = 8'h34;
        i_im2 = 8'h3A;
        i_im3 = 8'h38;
        i_im4 = 8'h32;
        i_im5 = 8'hB9;
        i_im6 = 8'hBC;
        i_im7 = 8'h3A;
        i_im8 = 8'h39;
        i_im9 = 8'h3A;
        #10 //15-15
        i_im1 = 8'h3A;
        i_im2 = 8'h38;
        i_im3 = 8'hB8;
        i_im4 = 8'hB9;
        i_im5 = 8'hBC;
        i_im6 = 8'hB9;
        i_im7 = 8'h39;
        i_im8 = 8'h3A;
        i_im9 = 8'h33;
        #10 //15-16
        i_im1 = 8'h38;
        i_im2 = 8'hB8;
        i_im3 = 8'hB1;
        i_im4 = 8'hBC;
        i_im5 = 8'hB9;
        i_im6 = 8'hBC;
        i_im7 = 8'h3A;
        i_im8 = 8'h33;
        i_im9 = 8'hAF;
        #10 //15-17
        i_im1 = 8'hB8;
        i_im2 = 8'hB1;
        i_im3 = 8'hB4;
        i_im4 = 8'hB9;
        i_im5 = 8'hBC;
        i_im6 = 8'hB4;
        i_im7 = 8'h33;
        i_im8 = 8'hAF;
        i_im9 = 8'h36;
        #10 //15-18
        i_im1 = 8'hB1;
        i_im2 = 8'hB4;
        i_im3 = 8'h32;
        i_im4 = 8'hBC;
        i_im5 = 8'hB4;
        i_im6 = 8'hA7;
        i_im7 = 8'hAF;
        i_im8 = 8'h36;
        i_im9 = 8'h39;
        #10 //15-19
        i_im1 = 8'hB4;
        i_im2 = 8'h32;
        i_im3 = 8'h37;
        i_im4 = 8'hB4;
        i_im5 = 8'hA7;
        i_im6 = 8'h20;
        i_im7 = 8'h36;
        i_im8 = 8'h39;
        i_im9 = 8'h2D;
        #10 //15-20
        i_im1 = 8'h32;
        i_im2 = 8'h37;
        i_im3 = 8'h3A;
        i_im4 = 8'hA7;
        i_im5 = 8'h20;
        i_im6 = 8'h28;
        i_im7 = 8'h39;
        i_im8 = 8'h2D;
        i_im9 = 8'hB9;
        #10 //15-21
        i_im1 = 8'h37;
        i_im2 = 8'h3A;
        i_im3 = 8'h2F;
        i_im4 = 8'h20;
        i_im5 = 8'h28;
        i_im6 = 8'hBA;
        i_im7 = 8'h2D;
        i_im8 = 8'hB9;
        i_im9 = 8'hB7;
        #10 //15-22
        i_im1 = 8'h3A;
        i_im2 = 8'h2F;
        i_im3 = 8'h3B;
        i_im4 = 8'h28;
        i_im5 = 8'hBA;
        i_im6 = 8'hBA;
        i_im7 = 8'hB9;
        i_im8 = 8'hB7;
        i_im9 = 8'hB0;
        #10 //15-23
        i_im1 = 8'h2F;
        i_im2 = 8'h3B;
        i_im3 = 8'h36;
        i_im4 = 8'hBA;
        i_im5 = 8'hBA;
        i_im6 = 8'h3A;
        i_im7 = 8'hB7;
        i_im8 = 8'hB0;
        i_im9 = 8'h38;
        #10 //15-24
        i_im1 = 8'h3B;
        i_im2 = 8'h36;
        i_im3 = 8'hBA;
        i_im4 = 8'hBA;
        i_im5 = 8'h3A;
        i_im6 = 8'h3B;
        i_im7 = 8'hB0;
        i_im8 = 8'h38;
        i_im9 = 8'h3B;
        #10 //15-25
        i_im1 = 8'h36;
        i_im2 = 8'hBA;
        i_im3 = 8'h3A;
        i_im4 = 8'h3A;
        i_im5 = 8'h3B;
        i_im6 = 8'h39;
        i_im7 = 8'h38;
        i_im8 = 8'h3B;
        i_im9 = 8'hB0;
        #10 //15-26
        i_im1 = 8'hBA;
        i_im2 = 8'h3A;
        i_im3 = 8'h34;
        i_im4 = 8'h3B;
        i_im5 = 8'h39;
        i_im6 = 8'hB9;
        i_im7 = 8'h3B;
        i_im8 = 8'hB0;
        i_im9 = 8'hB9;
        #10 //16-1
        i_im1 = 8'h2B;
        i_im2 = 8'h3C;
        i_im3 = 8'h2F;
        i_im4 = 8'h39;
        i_im5 = 8'h36;
        i_im6 = 8'hB3;
        i_im7 = 8'h3A;
        i_im8 = 8'hB6;
        i_im9 = 8'hBB;
        #10 //16-2
        i_im1 = 8'h3C;
        i_im2 = 8'h2F;
        i_im3 = 8'h3A;
        i_im4 = 8'h36;
        i_im5 = 8'hB3;
        i_im6 = 8'hB3;
        i_im7 = 8'hB6;
        i_im8 = 8'hBB;
        i_im9 = 8'h36;
        #10 //16-3
        i_im1 = 8'h2F;
        i_im2 = 8'h3A;
        i_im3 = 8'hB5;
        i_im4 = 8'hB3;
        i_im5 = 8'hB3;
        i_im6 = 8'hBA;
        i_im7 = 8'hBB;
        i_im8 = 8'h36;
        i_im9 = 8'hBA;
        #10 //16-4
        i_im1 = 8'h3A;
        i_im2 = 8'hB5;
        i_im3 = 8'h31;
        i_im4 = 8'hB3;
        i_im5 = 8'hBA;
        i_im6 = 8'hB9;
        i_im7 = 8'h36;
        i_im8 = 8'hBA;
        i_im9 = 8'hB5;
        #10 //16-5
        i_im1 = 8'hB5;
        i_im2 = 8'h31;
        i_im3 = 8'hB9;
        i_im4 = 8'hBA;
        i_im5 = 8'hB9;
        i_im6 = 8'hB5;
        i_im7 = 8'hBA;
        i_im8 = 8'hB5;
        i_im9 = 8'hB9;
        #10 //16-6
        i_im1 = 8'h31;
        i_im2 = 8'hB9;
        i_im3 = 8'h2B;
        i_im4 = 8'hB9;
        i_im5 = 8'hB5;
        i_im6 = 8'h3A;
        i_im7 = 8'hB5;
        i_im8 = 8'hB9;
        i_im9 = 8'hBB;
        #10 //16-7
        i_im1 = 8'hB9;
        i_im2 = 8'h2B;
        i_im3 = 8'hB2;
        i_im4 = 8'hB5;
        i_im5 = 8'h3A;
        i_im6 = 8'h2E;
        i_im7 = 8'hB9;
        i_im8 = 8'hBB;
        i_im9 = 8'hBB;
        #10 //16-8
        i_im1 = 8'h2B;
        i_im2 = 8'hB2;
        i_im3 = 8'hB9;
        i_im4 = 8'h3A;
        i_im5 = 8'h2E;
        i_im6 = 8'hB9;
        i_im7 = 8'hBB;
        i_im8 = 8'hBB;
        i_im9 = 8'hA9;
        #10 //16-9
        i_im1 = 8'hB2;
        i_im2 = 8'hB9;
        i_im3 = 8'hB5;
        i_im4 = 8'h2E;
        i_im5 = 8'hB9;
        i_im6 = 8'hBA;
        i_im7 = 8'hBB;
        i_im8 = 8'hA9;
        i_im9 = 8'hB9;
        #10 //16-10
        i_im1 = 8'hB9;
        i_im2 = 8'hB5;
        i_im3 = 8'hB8;
        i_im4 = 8'hB9;
        i_im5 = 8'hBA;
        i_im6 = 8'hB8;
        i_im7 = 8'hA9;
        i_im8 = 8'hB9;
        i_im9 = 8'h1C;
        #10 //16-11
        i_im1 = 8'hB5;
        i_im2 = 8'hB8;
        i_im3 = 8'hBA;
        i_im4 = 8'hBA;
        i_im5 = 8'hB8;
        i_im6 = 8'h35;
        i_im7 = 8'hB9;
        i_im8 = 8'h1C;
        i_im9 = 8'h37;
        #10 //16-12
        i_im1 = 8'hB8;
        i_im2 = 8'hBA;
        i_im3 = 8'h32;
        i_im4 = 8'hB8;
        i_im5 = 8'h35;
        i_im6 = 8'h3A;
        i_im7 = 8'h1C;
        i_im8 = 8'h37;
        i_im9 = 8'h32;
        #10 //16-13
        i_im1 = 8'hBA;
        i_im2 = 8'h32;
        i_im3 = 8'hB9;
        i_im4 = 8'h35;
        i_im5 = 8'h3A;
        i_im6 = 8'h39;
        i_im7 = 8'h37;
        i_im8 = 8'h32;
        i_im9 = 8'hBA;
        #10 //16-14
        i_im1 = 8'h32;
        i_im2 = 8'hB9;
        i_im3 = 8'hBC;
        i_im4 = 8'h3A;
        i_im5 = 8'h39;
        i_im6 = 8'h3A;
        i_im7 = 8'h32;
        i_im8 = 8'hBA;
        i_im9 = 8'h34;
        #10 //16-15
        i_im1 = 8'hB9;
        i_im2 = 8'hBC;
        i_im3 = 8'hB9;
        i_im4 = 8'h39;
        i_im5 = 8'h3A;
        i_im6 = 8'h33;
        i_im7 = 8'hBA;
        i_im8 = 8'h34;
        i_im9 = 8'hB7;
        #10 //16-16
        i_im1 = 8'hBC;
        i_im2 = 8'hB9;
        i_im3 = 8'hBC;
        i_im4 = 8'h3A;
        i_im5 = 8'h33;
        i_im6 = 8'hAF;
        i_im7 = 8'h34;
        i_im8 = 8'hB7;
        i_im9 = 8'hB0;
        #10 //16-17
        i_im1 = 8'hB9;
        i_im2 = 8'hBC;
        i_im3 = 8'hB4;
        i_im4 = 8'h33;
        i_im5 = 8'hAF;
        i_im6 = 8'h36;
        i_im7 = 8'hB7;
        i_im8 = 8'hB0;
        i_im9 = 8'hB2;
        #10 //16-18
        i_im1 = 8'hBC;
        i_im2 = 8'hB4;
        i_im3 = 8'hA7;
        i_im4 = 8'hAF;
        i_im5 = 8'h36;
        i_im6 = 8'h39;
        i_im7 = 8'hB0;
        i_im8 = 8'hB2;
        i_im9 = 8'hBB;
        #10 //16-19
        i_im1 = 8'hB4;
        i_im2 = 8'hA7;
        i_im3 = 8'h20;
        i_im4 = 8'h36;
        i_im5 = 8'h39;
        i_im6 = 8'h2D;
        i_im7 = 8'hB2;
        i_im8 = 8'hBB;
        i_im9 = 8'h32;
        #10 //16-20
        i_im1 = 8'hA7;
        i_im2 = 8'h20;
        i_im3 = 8'h28;
        i_im4 = 8'h39;
        i_im5 = 8'h2D;
        i_im6 = 8'hB9;
        i_im7 = 8'hBB;
        i_im8 = 8'h32;
        i_im9 = 8'h3B;
        #10 //16-21
        i_im1 = 8'h20;
        i_im2 = 8'h28;
        i_im3 = 8'hBA;
        i_im4 = 8'h2D;
        i_im5 = 8'hB9;
        i_im6 = 8'hB7;
        i_im7 = 8'h32;
        i_im8 = 8'h3B;
        i_im9 = 8'h2F;
        #10 //16-22
        i_im1 = 8'h28;
        i_im2 = 8'hBA;
        i_im3 = 8'hBA;
        i_im4 = 8'hB9;
        i_im5 = 8'hB7;
        i_im6 = 8'hB0;
        i_im7 = 8'h3B;
        i_im8 = 8'h2F;
        i_im9 = 8'h36;
        #10 //16-23
        i_im1 = 8'hBA;
        i_im2 = 8'hBA;
        i_im3 = 8'h3A;
        i_im4 = 8'hB7;
        i_im5 = 8'hB0;
        i_im6 = 8'h38;
        i_im7 = 8'h2F;
        i_im8 = 8'h36;
        i_im9 = 8'hB9;
        #10 //16-24
        i_im1 = 8'hBA;
        i_im2 = 8'h3A;
        i_im3 = 8'h3B;
        i_im4 = 8'hB0;
        i_im5 = 8'h38;
        i_im6 = 8'h3B;
        i_im7 = 8'h36;
        i_im8 = 8'hB9;
        i_im9 = 8'h31;
        #10 //16-25
        i_im1 = 8'h3A;
        i_im2 = 8'h3B;
        i_im3 = 8'h39;
        i_im4 = 8'h38;
        i_im5 = 8'h3B;
        i_im6 = 8'hB0;
        i_im7 = 8'hB9;
        i_im8 = 8'h31;
        i_im9 = 8'hAF;
        #10 //16-26
        i_im1 = 8'h3B;
        i_im2 = 8'h39;
        i_im3 = 8'hB9;
        i_im4 = 8'h3B;
        i_im5 = 8'hB0;
        i_im6 = 8'hB9;
        i_im7 = 8'h31;
        i_im8 = 8'hAF;
        i_im9 = 8'hBB;
        #10 //17-1
        i_im1 = 8'h39;
        i_im2 = 8'h36;
        i_im3 = 8'hB3;
        i_im4 = 8'h3A;
        i_im5 = 8'hB6;
        i_im6 = 8'hBB;
        i_im7 = 8'hB9;
        i_im8 = 8'hAC;
        i_im9 = 8'hB5;
        #10 //17-2
        i_im1 = 8'h36;
        i_im2 = 8'hB3;
        i_im3 = 8'hB3;
        i_im4 = 8'hB6;
        i_im5 = 8'hBB;
        i_im6 = 8'h36;
        i_im7 = 8'hAC;
        i_im8 = 8'hB5;
        i_im9 = 8'h3A;
        #10 //17-3
        i_im1 = 8'hB3;
        i_im2 = 8'hB3;
        i_im3 = 8'hBA;
        i_im4 = 8'hBB;
        i_im5 = 8'h36;
        i_im6 = 8'hBA;
        i_im7 = 8'hB5;
        i_im8 = 8'h3A;
        i_im9 = 8'hB5;
        #10 //17-4
        i_im1 = 8'hB3;
        i_im2 = 8'hBA;
        i_im3 = 8'hB9;
        i_im4 = 8'h36;
        i_im5 = 8'hBA;
        i_im6 = 8'hB5;
        i_im7 = 8'h3A;
        i_im8 = 8'hB5;
        i_im9 = 8'h37;
        #10 //17-5
        i_im1 = 8'hBA;
        i_im2 = 8'hB9;
        i_im3 = 8'hB5;
        i_im4 = 8'hBA;
        i_im5 = 8'hB5;
        i_im6 = 8'hB9;
        i_im7 = 8'hB5;
        i_im8 = 8'h37;
        i_im9 = 8'hB4;
        #10 //17-6
        i_im1 = 8'hB9;
        i_im2 = 8'hB5;
        i_im3 = 8'h3A;
        i_im4 = 8'hB5;
        i_im5 = 8'hB9;
        i_im6 = 8'hBB;
        i_im7 = 8'h37;
        i_im8 = 8'hB4;
        i_im9 = 8'hBC;
        #10 //17-7
        i_im1 = 8'hB5;
        i_im2 = 8'h3A;
        i_im3 = 8'h2E;
        i_im4 = 8'hB9;
        i_im5 = 8'hBB;
        i_im6 = 8'hBB;
        i_im7 = 8'hB4;
        i_im8 = 8'hBC;
        i_im9 = 8'h3B;
        #10 //17-8
        i_im1 = 8'h3A;
        i_im2 = 8'h2E;
        i_im3 = 8'hB9;
        i_im4 = 8'hBB;
        i_im5 = 8'hBB;
        i_im6 = 8'hA9;
        i_im7 = 8'hBC;
        i_im8 = 8'h3B;
        i_im9 = 8'hBB;
        #10 //17-9
        i_im1 = 8'h2E;
        i_im2 = 8'hB9;
        i_im3 = 8'hBA;
        i_im4 = 8'hBB;
        i_im5 = 8'hA9;
        i_im6 = 8'hB9;
        i_im7 = 8'h3B;
        i_im8 = 8'hBB;
        i_im9 = 8'hBC;
        #10 //17-10
        i_im1 = 8'hB9;
        i_im2 = 8'hBA;
        i_im3 = 8'hB8;
        i_im4 = 8'hA9;
        i_im5 = 8'hB9;
        i_im6 = 8'h1C;
        i_im7 = 8'hBB;
        i_im8 = 8'hBC;
        i_im9 = 8'hB9;
        #10 //17-11
        i_im1 = 8'hBA;
        i_im2 = 8'hB8;
        i_im3 = 8'h35;
        i_im4 = 8'hB9;
        i_im5 = 8'h1C;
        i_im6 = 8'h37;
        i_im7 = 8'hBC;
        i_im8 = 8'hB9;
        i_im9 = 8'hB4;
        #10 //17-12
        i_im1 = 8'hB8;
        i_im2 = 8'h35;
        i_im3 = 8'h3A;
        i_im4 = 8'h1C;
        i_im5 = 8'h37;
        i_im6 = 8'h32;
        i_im7 = 8'hB9;
        i_im8 = 8'hB4;
        i_im9 = 8'hBB;
        #10 //17-13
        i_im1 = 8'h35;
        i_im2 = 8'h3A;
        i_im3 = 8'h39;
        i_im4 = 8'h37;
        i_im5 = 8'h32;
        i_im6 = 8'hBA;
        i_im7 = 8'hB4;
        i_im8 = 8'hBB;
        i_im9 = 8'hB9;
        #10 //17-14
        i_im1 = 8'h3A;
        i_im2 = 8'h39;
        i_im3 = 8'h3A;
        i_im4 = 8'h32;
        i_im5 = 8'hBA;
        i_im6 = 8'h34;
        i_im7 = 8'hBB;
        i_im8 = 8'hB9;
        i_im9 = 8'h37;
        #10 //17-15
        i_im1 = 8'h39;
        i_im2 = 8'h3A;
        i_im3 = 8'h33;
        i_im4 = 8'hBA;
        i_im5 = 8'h34;
        i_im6 = 8'hB7;
        i_im7 = 8'hB9;
        i_im8 = 8'h37;
        i_im9 = 8'hB5;
        #10 //17-16
        i_im1 = 8'h3A;
        i_im2 = 8'h33;
        i_im3 = 8'hAF;
        i_im4 = 8'h34;
        i_im5 = 8'hB7;
        i_im6 = 8'hB0;
        i_im7 = 8'h37;
        i_im8 = 8'hB5;
        i_im9 = 8'h3B;
        #10 //17-17
        i_im1 = 8'h33;
        i_im2 = 8'hAF;
        i_im3 = 8'h36;
        i_im4 = 8'hB7;
        i_im5 = 8'hB0;
        i_im6 = 8'hB2;
        i_im7 = 8'hB5;
        i_im8 = 8'h3B;
        i_im9 = 8'h37;
        #10 //17-18
        i_im1 = 8'hAF;
        i_im2 = 8'h36;
        i_im3 = 8'h39;
        i_im4 = 8'hB0;
        i_im5 = 8'hB2;
        i_im6 = 8'hBB;
        i_im7 = 8'h3B;
        i_im8 = 8'h37;
        i_im9 = 8'hBA;
        #10 //17-19
        i_im1 = 8'h36;
        i_im2 = 8'h39;
        i_im3 = 8'h2D;
        i_im4 = 8'hB2;
        i_im5 = 8'hBB;
        i_im6 = 8'h32;
        i_im7 = 8'h37;
        i_im8 = 8'hBA;
        i_im9 = 8'hBB;
        #10 //17-20
        i_im1 = 8'h39;
        i_im2 = 8'h2D;
        i_im3 = 8'hB9;
        i_im4 = 8'hBB;
        i_im5 = 8'h32;
        i_im6 = 8'h3B;
        i_im7 = 8'hBA;
        i_im8 = 8'hBB;
        i_im9 = 8'h37;
        #10 //17-21
        i_im1 = 8'h2D;
        i_im2 = 8'hB9;
        i_im3 = 8'hB7;
        i_im4 = 8'h32;
        i_im5 = 8'h3B;
        i_im6 = 8'h2F;
        i_im7 = 8'hBB;
        i_im8 = 8'h37;
        i_im9 = 8'hBB;
        #10 //17-22
        i_im1 = 8'hB9;
        i_im2 = 8'hB7;
        i_im3 = 8'hB0;
        i_im4 = 8'h3B;
        i_im5 = 8'h2F;
        i_im6 = 8'h36;
        i_im7 = 8'h37;
        i_im8 = 8'hBB;
        i_im9 = 8'h30;
        #10 //17-23
        i_im1 = 8'hB7;
        i_im2 = 8'hB0;
        i_im3 = 8'h38;
        i_im4 = 8'h2F;
        i_im5 = 8'h36;
        i_im6 = 8'hB9;
        i_im7 = 8'hBB;
        i_im8 = 8'h30;
        i_im9 = 8'h26;
        #10 //17-24
        i_im1 = 8'hB0;
        i_im2 = 8'h38;
        i_im3 = 8'h3B;
        i_im4 = 8'h36;
        i_im5 = 8'hB9;
        i_im6 = 8'h31;
        i_im7 = 8'h30;
        i_im8 = 8'h26;
        i_im9 = 8'h3C;
        #10 //17-25
        i_im1 = 8'h38;
        i_im2 = 8'h3B;
        i_im3 = 8'hB0;
        i_im4 = 8'hB9;
        i_im5 = 8'h31;
        i_im6 = 8'hAF;
        i_im7 = 8'h26;
        i_im8 = 8'h3C;
        i_im9 = 8'hB5;
        #10 //17-26
        i_im1 = 8'h3B;
        i_im2 = 8'hB0;
        i_im3 = 8'hB9;
        i_im4 = 8'h31;
        i_im5 = 8'hAF;
        i_im6 = 8'hBB;
        i_im7 = 8'h3C;
        i_im8 = 8'hB5;
        i_im9 = 8'h39;
        #10 //18-1
        i_im1 = 8'h3A;
        i_im2 = 8'hB6;
        i_im3 = 8'hBB;
        i_im4 = 8'hB9;
        i_im5 = 8'hAC;
        i_im6 = 8'hB5;
        i_im7 = 8'h37;
        i_im8 = 8'hB2;
        i_im9 = 8'h32;
        #10 //18-2
        i_im1 = 8'hB6;
        i_im2 = 8'hBB;
        i_im3 = 8'h36;
        i_im4 = 8'hAC;
        i_im5 = 8'hB5;
        i_im6 = 8'h3A;
        i_im7 = 8'hB2;
        i_im8 = 8'h32;
        i_im9 = 8'h2F;
        #10 //18-3
        i_im1 = 8'hBB;
        i_im2 = 8'h36;
        i_im3 = 8'hBA;
        i_im4 = 8'hB5;
        i_im5 = 8'h3A;
        i_im6 = 8'hB5;
        i_im7 = 8'h32;
        i_im8 = 8'h2F;
        i_im9 = 8'hB3;
        #10 //18-4
        i_im1 = 8'h36;
        i_im2 = 8'hBA;
        i_im3 = 8'hB5;
        i_im4 = 8'h3A;
        i_im5 = 8'hB5;
        i_im6 = 8'h37;
        i_im7 = 8'h2F;
        i_im8 = 8'hB3;
        i_im9 = 8'hBA;
        #10 //18-5
        i_im1 = 8'hBA;
        i_im2 = 8'hB5;
        i_im3 = 8'hB9;
        i_im4 = 8'hB5;
        i_im5 = 8'h37;
        i_im6 = 8'hB4;
        i_im7 = 8'hB3;
        i_im8 = 8'hBA;
        i_im9 = 8'hAC;
        #10 //18-6
        i_im1 = 8'hB5;
        i_im2 = 8'hB9;
        i_im3 = 8'hBB;
        i_im4 = 8'h37;
        i_im5 = 8'hB4;
        i_im6 = 8'hBC;
        i_im7 = 8'hBA;
        i_im8 = 8'hAC;
        i_im9 = 8'h2D;
        #10 //18-7
        i_im1 = 8'hB9;
        i_im2 = 8'hBB;
        i_im3 = 8'hBB;
        i_im4 = 8'hB4;
        i_im5 = 8'hBC;
        i_im6 = 8'h3B;
        i_im7 = 8'hAC;
        i_im8 = 8'h2D;
        i_im9 = 8'h3B;
        #10 //18-8
        i_im1 = 8'hBB;
        i_im2 = 8'hBB;
        i_im3 = 8'hA9;
        i_im4 = 8'hBC;
        i_im5 = 8'h3B;
        i_im6 = 8'hBB;
        i_im7 = 8'h2D;
        i_im8 = 8'h3B;
        i_im9 = 8'hB9;
        #10 //18-9
        i_im1 = 8'hBB;
        i_im2 = 8'hA9;
        i_im3 = 8'hB9;
        i_im4 = 8'h3B;
        i_im5 = 8'hBB;
        i_im6 = 8'hBC;
        i_im7 = 8'h3B;
        i_im8 = 8'hB9;
        i_im9 = 8'h36;
        #10 //18-10
        i_im1 = 8'hA9;
        i_im2 = 8'hB9;
        i_im3 = 8'h1C;
        i_im4 = 8'hBB;
        i_im5 = 8'hBC;
        i_im6 = 8'hB9;
        i_im7 = 8'hB9;
        i_im8 = 8'h36;
        i_im9 = 8'hAF;
        #10 //18-11
        i_im1 = 8'hB9;
        i_im2 = 8'h1C;
        i_im3 = 8'h37;
        i_im4 = 8'hBC;
        i_im5 = 8'hB9;
        i_im6 = 8'hB4;
        i_im7 = 8'h36;
        i_im8 = 8'hAF;
        i_im9 = 8'hBB;
        #10 //18-12
        i_im1 = 8'h1C;
        i_im2 = 8'h37;
        i_im3 = 8'h32;
        i_im4 = 8'hB9;
        i_im5 = 8'hB4;
        i_im6 = 8'hBB;
        i_im7 = 8'hAF;
        i_im8 = 8'hBB;
        i_im9 = 8'hB8;
        #10 //18-13
        i_im1 = 8'h37;
        i_im2 = 8'h32;
        i_im3 = 8'hBA;
        i_im4 = 8'hB4;
        i_im5 = 8'hBB;
        i_im6 = 8'hB9;
        i_im7 = 8'hBB;
        i_im8 = 8'hB8;
        i_im9 = 8'h35;
        #10 //18-14
        i_im1 = 8'h32;
        i_im2 = 8'hBA;
        i_im3 = 8'h34;
        i_im4 = 8'hBB;
        i_im5 = 8'hB9;
        i_im6 = 8'h37;
        i_im7 = 8'hB8;
        i_im8 = 8'h35;
        i_im9 = 8'h38;
        #10 //18-15
        i_im1 = 8'hBA;
        i_im2 = 8'h34;
        i_im3 = 8'hB7;
        i_im4 = 8'hB9;
        i_im5 = 8'h37;
        i_im6 = 8'hB5;
        i_im7 = 8'h35;
        i_im8 = 8'h38;
        i_im9 = 8'hB6;
        #10 //18-16
        i_im1 = 8'h34;
        i_im2 = 8'hB7;
        i_im3 = 8'hB0;
        i_im4 = 8'h37;
        i_im5 = 8'hB5;
        i_im6 = 8'h3B;
        i_im7 = 8'h38;
        i_im8 = 8'hB6;
        i_im9 = 8'h3C;
        #10 //18-17
        i_im1 = 8'hB7;
        i_im2 = 8'hB0;
        i_im3 = 8'hB2;
        i_im4 = 8'hB5;
        i_im5 = 8'h3B;
        i_im6 = 8'h37;
        i_im7 = 8'hB6;
        i_im8 = 8'h3C;
        i_im9 = 8'hB3;
        #10 //18-18
        i_im1 = 8'hB0;
        i_im2 = 8'hB2;
        i_im3 = 8'hBB;
        i_im4 = 8'h3B;
        i_im5 = 8'h37;
        i_im6 = 8'hBA;
        i_im7 = 8'h3C;
        i_im8 = 8'hB3;
        i_im9 = 8'h3B;
        #10 //18-19
        i_im1 = 8'hB2;
        i_im2 = 8'hBB;
        i_im3 = 8'h32;
        i_im4 = 8'h37;
        i_im5 = 8'hBA;
        i_im6 = 8'hBB;
        i_im7 = 8'hB3;
        i_im8 = 8'h3B;
        i_im9 = 8'hBB;
        #10 //18-20
        i_im1 = 8'hBB;
        i_im2 = 8'h32;
        i_im3 = 8'h3B;
        i_im4 = 8'hBA;
        i_im5 = 8'hBB;
        i_im6 = 8'h37;
        i_im7 = 8'h3B;
        i_im8 = 8'hBB;
        i_im9 = 8'hB6;
        #10 //18-21
        i_im1 = 8'h32;
        i_im2 = 8'h3B;
        i_im3 = 8'h2F;
        i_im4 = 8'hBB;
        i_im5 = 8'h37;
        i_im6 = 8'hBB;
        i_im7 = 8'hBB;
        i_im8 = 8'hB6;
        i_im9 = 8'hB3;
        #10 //18-22
        i_im1 = 8'h3B;
        i_im2 = 8'h2F;
        i_im3 = 8'h36;
        i_im4 = 8'h37;
        i_im5 = 8'hBB;
        i_im6 = 8'h30;
        i_im7 = 8'hB6;
        i_im8 = 8'hB3;
        i_im9 = 8'hBB;
        #10 //18-23
        i_im1 = 8'h2F;
        i_im2 = 8'h36;
        i_im3 = 8'hB9;
        i_im4 = 8'hBB;
        i_im5 = 8'h30;
        i_im6 = 8'h26;
        i_im7 = 8'hB3;
        i_im8 = 8'hBB;
        i_im9 = 8'hBB;
        #10 //18-24
        i_im1 = 8'h36;
        i_im2 = 8'hB9;
        i_im3 = 8'h31;
        i_im4 = 8'h30;
        i_im5 = 8'h26;
        i_im6 = 8'h3C;
        i_im7 = 8'hBB;
        i_im8 = 8'hBB;
        i_im9 = 8'h37;
        #10 //18-25
        i_im1 = 8'hB9;
        i_im2 = 8'h31;
        i_im3 = 8'hAF;
        i_im4 = 8'h26;
        i_im5 = 8'h3C;
        i_im6 = 8'hB5;
        i_im7 = 8'hBB;
        i_im8 = 8'h37;
        i_im9 = 8'hB3;
        #10 //18-26
        i_im1 = 8'h31;
        i_im2 = 8'hAF;
        i_im3 = 8'hBB;
        i_im4 = 8'h3C;
        i_im5 = 8'hB5;
        i_im6 = 8'h39;
        i_im7 = 8'h37;
        i_im8 = 8'hB3;
        i_im9 = 8'hBB;
        #10 //19-1
        i_im1 = 8'hB9;
        i_im2 = 8'hAC;
        i_im3 = 8'hB5;
        i_im4 = 8'h37;
        i_im5 = 8'hB2;
        i_im6 = 8'h32;
        i_im7 = 8'hBB;
        i_im8 = 8'hB4;
        i_im9 = 8'hB4;
        #10 //19-2
        i_im1 = 8'hAC;
        i_im2 = 8'hB5;
        i_im3 = 8'h3A;
        i_im4 = 8'hB2;
        i_im5 = 8'h32;
        i_im6 = 8'h2F;
        i_im7 = 8'hB4;
        i_im8 = 8'hB4;
        i_im9 = 8'h37;
        #10 //19-3
        i_im1 = 8'hB5;
        i_im2 = 8'h3A;
        i_im3 = 8'hB5;
        i_im4 = 8'h32;
        i_im5 = 8'h2F;
        i_im6 = 8'hB3;
        i_im7 = 8'hB4;
        i_im8 = 8'h37;
        i_im9 = 8'hB7;
        #10 //19-4
        i_im1 = 8'h3A;
        i_im2 = 8'hB5;
        i_im3 = 8'h37;
        i_im4 = 8'h2F;
        i_im5 = 8'hB3;
        i_im6 = 8'hBA;
        i_im7 = 8'h37;
        i_im8 = 8'hB7;
        i_im9 = 8'h3B;
        #10 //19-5
        i_im1 = 8'hB5;
        i_im2 = 8'h37;
        i_im3 = 8'hB4;
        i_im4 = 8'hB3;
        i_im5 = 8'hBA;
        i_im6 = 8'hAC;
        i_im7 = 8'hB7;
        i_im8 = 8'h3B;
        i_im9 = 8'h20;
        #10 //19-6
        i_im1 = 8'h37;
        i_im2 = 8'hB4;
        i_im3 = 8'hBC;
        i_im4 = 8'hBA;
        i_im5 = 8'hAC;
        i_im6 = 8'h2D;
        i_im7 = 8'h3B;
        i_im8 = 8'h20;
        i_im9 = 8'hBB;
        #10 //19-7
        i_im1 = 8'hB4;
        i_im2 = 8'hBC;
        i_im3 = 8'h3B;
        i_im4 = 8'hAC;
        i_im5 = 8'h2D;
        i_im6 = 8'h3B;
        i_im7 = 8'h20;
        i_im8 = 8'hBB;
        i_im9 = 8'hB9;
        #10 //19-8
        i_im1 = 8'hBC;
        i_im2 = 8'h3B;
        i_im3 = 8'hBB;
        i_im4 = 8'h2D;
        i_im5 = 8'h3B;
        i_im6 = 8'hB9;
        i_im7 = 8'hBB;
        i_im8 = 8'hB9;
        i_im9 = 8'h2E;
        #10 //19-9
        i_im1 = 8'h3B;
        i_im2 = 8'hBB;
        i_im3 = 8'hBC;
        i_im4 = 8'h3B;
        i_im5 = 8'hB9;
        i_im6 = 8'h36;
        i_im7 = 8'hB9;
        i_im8 = 8'h2E;
        i_im9 = 8'h2C;
        #10 //19-10
        i_im1 = 8'hBB;
        i_im2 = 8'hBC;
        i_im3 = 8'hB9;
        i_im4 = 8'hB9;
        i_im5 = 8'h36;
        i_im6 = 8'hAF;
        i_im7 = 8'h2E;
        i_im8 = 8'h2C;
        i_im9 = 8'hBA;
        #10 //19-11
        i_im1 = 8'hBC;
        i_im2 = 8'hB9;
        i_im3 = 8'hB4;
        i_im4 = 8'h36;
        i_im5 = 8'hAF;
        i_im6 = 8'hBB;
        i_im7 = 8'h2C;
        i_im8 = 8'hBA;
        i_im9 = 8'hBB;
        #10 //19-12
        i_im1 = 8'hB9;
        i_im2 = 8'hB4;
        i_im3 = 8'hBB;
        i_im4 = 8'hAF;
        i_im5 = 8'hBB;
        i_im6 = 8'hB8;
        i_im7 = 8'hBA;
        i_im8 = 8'hBB;
        i_im9 = 8'hBB;
        #10 //19-13
        i_im1 = 8'hB4;
        i_im2 = 8'hBB;
        i_im3 = 8'hB9;
        i_im4 = 8'hBB;
        i_im5 = 8'hB8;
        i_im6 = 8'h35;
        i_im7 = 8'hBB;
        i_im8 = 8'hBB;
        i_im9 = 8'h3B;
        #10 //19-14
        i_im1 = 8'hBB;
        i_im2 = 8'hB9;
        i_im3 = 8'h37;
        i_im4 = 8'hB8;
        i_im5 = 8'h35;
        i_im6 = 8'h38;
        i_im7 = 8'hBB;
        i_im8 = 8'h3B;
        i_im9 = 8'hBB;
        #10 //19-15
        i_im1 = 8'hB9;
        i_im2 = 8'h37;
        i_im3 = 8'hB5;
        i_im4 = 8'h35;
        i_im5 = 8'h38;
        i_im6 = 8'hB6;
        i_im7 = 8'h3B;
        i_im8 = 8'hBB;
        i_im9 = 8'hA5;
        #10 //19-16
        i_im1 = 8'h37;
        i_im2 = 8'hB5;
        i_im3 = 8'h3B;
        i_im4 = 8'h38;
        i_im5 = 8'hB6;
        i_im6 = 8'h3C;
        i_im7 = 8'hBB;
        i_im8 = 8'hA5;
        i_im9 = 8'h31;
        #10 //19-17
        i_im1 = 8'hB5;
        i_im2 = 8'h3B;
        i_im3 = 8'h37;
        i_im4 = 8'hB6;
        i_im5 = 8'h3C;
        i_im6 = 8'hB3;
        i_im7 = 8'hA5;
        i_im8 = 8'h31;
        i_im9 = 8'h39;
        #10 //19-18
        i_im1 = 8'h3B;
        i_im2 = 8'h37;
        i_im3 = 8'hBA;
        i_im4 = 8'h3C;
        i_im5 = 8'hB3;
        i_im6 = 8'h3B;
        i_im7 = 8'h31;
        i_im8 = 8'h39;
        i_im9 = 8'h35;
        #10 //19-19
        i_im1 = 8'h37;
        i_im2 = 8'hBA;
        i_im3 = 8'hBB;
        i_im4 = 8'hB3;
        i_im5 = 8'h3B;
        i_im6 = 8'hBB;
        i_im7 = 8'h39;
        i_im8 = 8'h35;
        i_im9 = 8'hB4;
        #10 //19-20
        i_im1 = 8'hBA;
        i_im2 = 8'hBB;
        i_im3 = 8'h37;
        i_im4 = 8'h3B;
        i_im5 = 8'hBB;
        i_im6 = 8'hB6;
        i_im7 = 8'h35;
        i_im8 = 8'hB4;
        i_im9 = 8'h38;
        #10 //19-21
        i_im1 = 8'hBB;
        i_im2 = 8'h37;
        i_im3 = 8'hBB;
        i_im4 = 8'hBB;
        i_im5 = 8'hB6;
        i_im6 = 8'hB3;
        i_im7 = 8'hB4;
        i_im8 = 8'h38;
        i_im9 = 8'hBA;
        #10 //19-22
        i_im1 = 8'h37;
        i_im2 = 8'hBB;
        i_im3 = 8'h30;
        i_im4 = 8'hB6;
        i_im5 = 8'hB3;
        i_im6 = 8'hBB;
        i_im7 = 8'h38;
        i_im8 = 8'hBA;
        i_im9 = 8'h37;
        #10 //19-23
        i_im1 = 8'hBB;
        i_im2 = 8'h30;
        i_im3 = 8'h26;
        i_im4 = 8'hB3;
        i_im5 = 8'hBB;
        i_im6 = 8'hBB;
        i_im7 = 8'hBA;
        i_im8 = 8'h37;
        i_im9 = 8'hB5;
        #10 //19-24
        i_im1 = 8'h30;
        i_im2 = 8'h26;
        i_im3 = 8'h3C;
        i_im4 = 8'hBB;
        i_im5 = 8'hBB;
        i_im6 = 8'h37;
        i_im7 = 8'h37;
        i_im8 = 8'hB5;
        i_im9 = 8'hB4;
        #10 //19-25
        i_im1 = 8'h26;
        i_im2 = 8'h3C;
        i_im3 = 8'hB5;
        i_im4 = 8'hBB;
        i_im5 = 8'h37;
        i_im6 = 8'hB3;
        i_im7 = 8'hB5;
        i_im8 = 8'hB4;
        i_im9 = 8'h2F;
        #10 //19-26
        i_im1 = 8'h3C;
        i_im2 = 8'hB5;
        i_im3 = 8'h39;
        i_im4 = 8'h37;
        i_im5 = 8'hB3;
        i_im6 = 8'hBB;
        i_im7 = 8'hB4;
        i_im8 = 8'h2F;
        i_im9 = 8'hB8;
        #10 //20-1
        i_im1 = 8'h37;
        i_im2 = 8'hB2;
        i_im3 = 8'h32;
        i_im4 = 8'hBB;
        i_im5 = 8'hB4;
        i_im6 = 8'hB4;
        i_im7 = 8'h3B;
        i_im8 = 8'hBA;
        i_im9 = 8'hAD;
        #10 //20-2
        i_im1 = 8'hB2;
        i_im2 = 8'h32;
        i_im3 = 8'h2F;
        i_im4 = 8'hB4;
        i_im5 = 8'hB4;
        i_im6 = 8'h37;
        i_im7 = 8'hBA;
        i_im8 = 8'hAD;
        i_im9 = 8'h3B;
        #10 //20-3
        i_im1 = 8'h32;
        i_im2 = 8'h2F;
        i_im3 = 8'hB3;
        i_im4 = 8'hB4;
        i_im5 = 8'h37;
        i_im6 = 8'hB7;
        i_im7 = 8'hAD;
        i_im8 = 8'h3B;
        i_im9 = 8'h3B;
        #10 //20-4
        i_im1 = 8'h2F;
        i_im2 = 8'hB3;
        i_im3 = 8'hBA;
        i_im4 = 8'h37;
        i_im5 = 8'hB7;
        i_im6 = 8'h3B;
        i_im7 = 8'h3B;
        i_im8 = 8'h3B;
        i_im9 = 8'h39;
        #10 //20-5
        i_im1 = 8'hB3;
        i_im2 = 8'hBA;
        i_im3 = 8'hAC;
        i_im4 = 8'hB7;
        i_im5 = 8'h3B;
        i_im6 = 8'h20;
        i_im7 = 8'h3B;
        i_im8 = 8'h39;
        i_im9 = 8'h37;
        #10 //20-6
        i_im1 = 8'hBA;
        i_im2 = 8'hAC;
        i_im3 = 8'h2D;
        i_im4 = 8'h3B;
        i_im5 = 8'h20;
        i_im6 = 8'hBB;
        i_im7 = 8'h39;
        i_im8 = 8'h37;
        i_im9 = 8'h3B;
        #10 //20-7
        i_im1 = 8'hAC;
        i_im2 = 8'h2D;
        i_im3 = 8'h3B;
        i_im4 = 8'h20;
        i_im5 = 8'hBB;
        i_im6 = 8'hB9;
        i_im7 = 8'h37;
        i_im8 = 8'h3B;
        i_im9 = 8'hB8;
        #10 //20-8
        i_im1 = 8'h2D;
        i_im2 = 8'h3B;
        i_im3 = 8'hB9;
        i_im4 = 8'hBB;
        i_im5 = 8'hB9;
        i_im6 = 8'h2E;
        i_im7 = 8'h3B;
        i_im8 = 8'hB8;
        i_im9 = 8'h39;
        #10 //20-9
        i_im1 = 8'h3B;
        i_im2 = 8'hB9;
        i_im3 = 8'h36;
        i_im4 = 8'hB9;
        i_im5 = 8'h2E;
        i_im6 = 8'h2C;
        i_im7 = 8'hB8;
        i_im8 = 8'h39;
        i_im9 = 8'hB6;
        #10 //20-10
        i_im1 = 8'hB9;
        i_im2 = 8'h36;
        i_im3 = 8'hAF;
        i_im4 = 8'h2E;
        i_im5 = 8'h2C;
        i_im6 = 8'hBA;
        i_im7 = 8'h39;
        i_im8 = 8'hB6;
        i_im9 = 8'hB6;
        #10 //20-11
        i_im1 = 8'h36;
        i_im2 = 8'hAF;
        i_im3 = 8'hBB;
        i_im4 = 8'h2C;
        i_im5 = 8'hBA;
        i_im6 = 8'hBB;
        i_im7 = 8'hB6;
        i_im8 = 8'hB6;
        i_im9 = 8'hA0;
        #10 //20-12
        i_im1 = 8'hAF;
        i_im2 = 8'hBB;
        i_im3 = 8'hB8;
        i_im4 = 8'hBA;
        i_im5 = 8'hBB;
        i_im6 = 8'hBB;
        i_im7 = 8'hB6;
        i_im8 = 8'hA0;
        i_im9 = 8'h38;
        #10 //20-13
        i_im1 = 8'hBB;
        i_im2 = 8'hB8;
        i_im3 = 8'h35;
        i_im4 = 8'hBB;
        i_im5 = 8'hBB;
        i_im6 = 8'h3B;
        i_im7 = 8'hA0;
        i_im8 = 8'h38;
        i_im9 = 8'h3B;
        #10 //20-14
        i_im1 = 8'hB8;
        i_im2 = 8'h35;
        i_im3 = 8'h38;
        i_im4 = 8'hBB;
        i_im5 = 8'h3B;
        i_im6 = 8'hBB;
        i_im7 = 8'h38;
        i_im8 = 8'h3B;
        i_im9 = 8'h38;
        #10 //20-15
        i_im1 = 8'h35;
        i_im2 = 8'h38;
        i_im3 = 8'hB6;
        i_im4 = 8'h3B;
        i_im5 = 8'hBB;
        i_im6 = 8'hA5;
        i_im7 = 8'h3B;
        i_im8 = 8'h38;
        i_im9 = 8'hBB;
        #10 //20-16
        i_im1 = 8'h38;
        i_im2 = 8'hB6;
        i_im3 = 8'h3C;
        i_im4 = 8'hBB;
        i_im5 = 8'hA5;
        i_im6 = 8'h31;
        i_im7 = 8'h38;
        i_im8 = 8'hBB;
        i_im9 = 8'h39;
        #10 //20-17
        i_im1 = 8'hB6;
        i_im2 = 8'h3C;
        i_im3 = 8'hB3;
        i_im4 = 8'hA5;
        i_im5 = 8'h31;
        i_im6 = 8'h39;
        i_im7 = 8'hBB;
        i_im8 = 8'h39;
        i_im9 = 8'h35;
        #10 //20-18
        i_im1 = 8'h3C;
        i_im2 = 8'hB3;
        i_im3 = 8'h3B;
        i_im4 = 8'h31;
        i_im5 = 8'h39;
        i_im6 = 8'h35;
        i_im7 = 8'h39;
        i_im8 = 8'h35;
        i_im9 = 8'hAF;
        #10 //20-19
        i_im1 = 8'hB3;
        i_im2 = 8'h3B;
        i_im3 = 8'hBB;
        i_im4 = 8'h39;
        i_im5 = 8'h35;
        i_im6 = 8'hB4;
        i_im7 = 8'h35;
        i_im8 = 8'hAF;
        i_im9 = 8'hB8;
        #10 //20-20
        i_im1 = 8'h3B;
        i_im2 = 8'hBB;
        i_im3 = 8'hB6;
        i_im4 = 8'h35;
        i_im5 = 8'hB4;
        i_im6 = 8'h38;
        i_im7 = 8'hAF;
        i_im8 = 8'hB8;
        i_im9 = 8'h38;
        #10 //20-21
        i_im1 = 8'hBB;
        i_im2 = 8'hB6;
        i_im3 = 8'hB3;
        i_im4 = 8'hB4;
        i_im5 = 8'h38;
        i_im6 = 8'hBA;
        i_im7 = 8'hB8;
        i_im8 = 8'h38;
        i_im9 = 8'h3A;
        #10 //20-22
        i_im1 = 8'hB6;
        i_im2 = 8'hB3;
        i_im3 = 8'hBB;
        i_im4 = 8'h38;
        i_im5 = 8'hBA;
        i_im6 = 8'h37;
        i_im7 = 8'h38;
        i_im8 = 8'h3A;
        i_im9 = 8'h38;
        #10 //20-23
        i_im1 = 8'hB3;
        i_im2 = 8'hBB;
        i_im3 = 8'hBB;
        i_im4 = 8'hBA;
        i_im5 = 8'h37;
        i_im6 = 8'hB5;
        i_im7 = 8'h3A;
        i_im8 = 8'h38;
        i_im9 = 8'hAE;
        #10 //20-24
        i_im1 = 8'hBB;
        i_im2 = 8'hBB;
        i_im3 = 8'h37;
        i_im4 = 8'h37;
        i_im5 = 8'hB5;
        i_im6 = 8'hB4;
        i_im7 = 8'h38;
        i_im8 = 8'hAE;
        i_im9 = 8'h34;
        #10 //20-25
        i_im1 = 8'hBB;
        i_im2 = 8'h37;
        i_im3 = 8'hB3;
        i_im4 = 8'hB5;
        i_im5 = 8'hB4;
        i_im6 = 8'h2F;
        i_im7 = 8'hAE;
        i_im8 = 8'h34;
        i_im9 = 8'h36;
        #10 //20-26
        i_im1 = 8'h37;
        i_im2 = 8'hB3;
        i_im3 = 8'hBB;
        i_im4 = 8'hB4;
        i_im5 = 8'h2F;
        i_im6 = 8'hB8;
        i_im7 = 8'h34;
        i_im8 = 8'h36;
        i_im9 = 8'h39;
        #10 //21-1
        i_im1 = 8'hBB;
        i_im2 = 8'hB4;
        i_im3 = 8'hB4;
        i_im4 = 8'h3B;
        i_im5 = 8'hBA;
        i_im6 = 8'hAD;
        i_im7 = 8'h39;
        i_im8 = 8'hB6;
        i_im9 = 8'hBA;
        #10 //21-2
        i_im1 = 8'hB4;
        i_im2 = 8'hB4;
        i_im3 = 8'h37;
        i_im4 = 8'hBA;
        i_im5 = 8'hAD;
        i_im6 = 8'h3B;
        i_im7 = 8'hB6;
        i_im8 = 8'hBA;
        i_im9 = 8'hB9;
        #10 //21-3
        i_im1 = 8'hB4;
        i_im2 = 8'h37;
        i_im3 = 8'hB7;
        i_im4 = 8'hAD;
        i_im5 = 8'h3B;
        i_im6 = 8'h3B;
        i_im7 = 8'hBA;
        i_im8 = 8'hB9;
        i_im9 = 8'h39;
        #10 //21-4
        i_im1 = 8'h37;
        i_im2 = 8'hB7;
        i_im3 = 8'h3B;
        i_im4 = 8'h3B;
        i_im5 = 8'h3B;
        i_im6 = 8'h39;
        i_im7 = 8'hB9;
        i_im8 = 8'h39;
        i_im9 = 8'h38;
        #10 //21-5
        i_im1 = 8'hB7;
        i_im2 = 8'h3B;
        i_im3 = 8'h20;
        i_im4 = 8'h3B;
        i_im5 = 8'h39;
        i_im6 = 8'h37;
        i_im7 = 8'h39;
        i_im8 = 8'h38;
        i_im9 = 8'hB5;
        #10 //21-6
        i_im1 = 8'h3B;
        i_im2 = 8'h20;
        i_im3 = 8'hBB;
        i_im4 = 8'h39;
        i_im5 = 8'h37;
        i_im6 = 8'h3B;
        i_im7 = 8'h38;
        i_im8 = 8'hB5;
        i_im9 = 8'hB6;
        #10 //21-7
        i_im1 = 8'h20;
        i_im2 = 8'hBB;
        i_im3 = 8'hB9;
        i_im4 = 8'h37;
        i_im5 = 8'h3B;
        i_im6 = 8'hB8;
        i_im7 = 8'hB5;
        i_im8 = 8'hB6;
        i_im9 = 8'hBB;
        #10 //21-8
        i_im1 = 8'hBB;
        i_im2 = 8'hB9;
        i_im3 = 8'h2E;
        i_im4 = 8'h3B;
        i_im5 = 8'hB8;
        i_im6 = 8'h39;
        i_im7 = 8'hB6;
        i_im8 = 8'hBB;
        i_im9 = 8'h3B;
        #10 //21-9
        i_im1 = 8'hB9;
        i_im2 = 8'h2E;
        i_im3 = 8'h2C;
        i_im4 = 8'hB8;
        i_im5 = 8'h39;
        i_im6 = 8'hB6;
        i_im7 = 8'hBB;
        i_im8 = 8'h3B;
        i_im9 = 8'h39;
        #10 //21-10
        i_im1 = 8'h2E;
        i_im2 = 8'h2C;
        i_im3 = 8'hBA;
        i_im4 = 8'h39;
        i_im5 = 8'hB6;
        i_im6 = 8'hB6;
        i_im7 = 8'h3B;
        i_im8 = 8'h39;
        i_im9 = 8'h3B;
        #10 //21-11
        i_im1 = 8'h2C;
        i_im2 = 8'hBA;
        i_im3 = 8'hBB;
        i_im4 = 8'hB6;
        i_im5 = 8'hB6;
        i_im6 = 8'hA0;
        i_im7 = 8'h39;
        i_im8 = 8'h3B;
        i_im9 = 8'hB0;
        #10 //21-12
        i_im1 = 8'hBA;
        i_im2 = 8'hBB;
        i_im3 = 8'hBB;
        i_im4 = 8'hB6;
        i_im5 = 8'hA0;
        i_im6 = 8'h38;
        i_im7 = 8'h3B;
        i_im8 = 8'hB0;
        i_im9 = 8'hBC;
        #10 //21-13
        i_im1 = 8'hBB;
        i_im2 = 8'hBB;
        i_im3 = 8'h3B;
        i_im4 = 8'hA0;
        i_im5 = 8'h38;
        i_im6 = 8'h3B;
        i_im7 = 8'hB0;
        i_im8 = 8'hBC;
        i_im9 = 8'hB5;
        #10 //21-14
        i_im1 = 8'hBB;
        i_im2 = 8'h3B;
        i_im3 = 8'hBB;
        i_im4 = 8'h38;
        i_im5 = 8'h3B;
        i_im6 = 8'h38;
        i_im7 = 8'hBC;
        i_im8 = 8'hB5;
        i_im9 = 8'hB4;
        #10 //21-15
        i_im1 = 8'h3B;
        i_im2 = 8'hBB;
        i_im3 = 8'hA5;
        i_im4 = 8'h3B;
        i_im5 = 8'h38;
        i_im6 = 8'hBB;
        i_im7 = 8'hB5;
        i_im8 = 8'hB4;
        i_im9 = 8'hB9;
        #10 //21-16
        i_im1 = 8'hBB;
        i_im2 = 8'hA5;
        i_im3 = 8'h31;
        i_im4 = 8'h38;
        i_im5 = 8'hBB;
        i_im6 = 8'h39;
        i_im7 = 8'hB4;
        i_im8 = 8'hB9;
        i_im9 = 8'h30;
        #10 //21-17
        i_im1 = 8'hA5;
        i_im2 = 8'h31;
        i_im3 = 8'h39;
        i_im4 = 8'hBB;
        i_im5 = 8'h39;
        i_im6 = 8'h35;
        i_im7 = 8'hB9;
        i_im8 = 8'h30;
        i_im9 = 8'hBA;
        #10 //21-18
        i_im1 = 8'h31;
        i_im2 = 8'h39;
        i_im3 = 8'h35;
        i_im4 = 8'h39;
        i_im5 = 8'h35;
        i_im6 = 8'hAF;
        i_im7 = 8'h30;
        i_im8 = 8'hBA;
        i_im9 = 8'h39;
        #10 //21-19
        i_im1 = 8'h39;
        i_im2 = 8'h35;
        i_im3 = 8'hB4;
        i_im4 = 8'h35;
        i_im5 = 8'hAF;
        i_im6 = 8'hB8;
        i_im7 = 8'hBA;
        i_im8 = 8'h39;
        i_im9 = 8'hB8;
        #10 //21-20
        i_im1 = 8'h35;
        i_im2 = 8'hB4;
        i_im3 = 8'h38;
        i_im4 = 8'hAF;
        i_im5 = 8'hB8;
        i_im6 = 8'h38;
        i_im7 = 8'h39;
        i_im8 = 8'hB8;
        i_im9 = 8'hBB;
        #10 //21-21
        i_im1 = 8'hB4;
        i_im2 = 8'h38;
        i_im3 = 8'hBA;
        i_im4 = 8'hB8;
        i_im5 = 8'h38;
        i_im6 = 8'h3A;
        i_im7 = 8'hB8;
        i_im8 = 8'hBB;
        i_im9 = 8'h3B;
        #10 //21-22
        i_im1 = 8'h38;
        i_im2 = 8'hBA;
        i_im3 = 8'h37;
        i_im4 = 8'h38;
        i_im5 = 8'h3A;
        i_im6 = 8'h38;
        i_im7 = 8'hBB;
        i_im8 = 8'h3B;
        i_im9 = 8'h35;
        #10 //21-23
        i_im1 = 8'hBA;
        i_im2 = 8'h37;
        i_im3 = 8'hB5;
        i_im4 = 8'h3A;
        i_im5 = 8'h38;
        i_im6 = 8'hAE;
        i_im7 = 8'h3B;
        i_im8 = 8'h35;
        i_im9 = 8'h3C;
        #10 //21-24
        i_im1 = 8'h37;
        i_im2 = 8'hB5;
        i_im3 = 8'hB4;
        i_im4 = 8'h38;
        i_im5 = 8'hAE;
        i_im6 = 8'h34;
        i_im7 = 8'h35;
        i_im8 = 8'h3C;
        i_im9 = 8'h39;
        #10 //21-25
        i_im1 = 8'hB5;
        i_im2 = 8'hB4;
        i_im3 = 8'h2F;
        i_im4 = 8'hAE;
        i_im5 = 8'h34;
        i_im6 = 8'h36;
        i_im7 = 8'h3C;
        i_im8 = 8'h39;
        i_im9 = 8'h3A;
        #10 //21-26
        i_im1 = 8'hB4;
        i_im2 = 8'h2F;
        i_im3 = 8'hB8;
        i_im4 = 8'h34;
        i_im5 = 8'h36;
        i_im6 = 8'h39;
        i_im7 = 8'h39;
        i_im8 = 8'h3A;
        i_im9 = 8'hB2;
        #10 //22-1
        i_im1 = 8'h3B;
        i_im2 = 8'hBA;
        i_im3 = 8'hAD;
        i_im4 = 8'h39;
        i_im5 = 8'hB6;
        i_im6 = 8'hBA;
        i_im7 = 8'hBA;
        i_im8 = 8'h36;
        i_im9 = 8'h37;
        #10 //22-2
        i_im1 = 8'hBA;
        i_im2 = 8'hAD;
        i_im3 = 8'h3B;
        i_im4 = 8'hB6;
        i_im5 = 8'hBA;
        i_im6 = 8'hB9;
        i_im7 = 8'h36;
        i_im8 = 8'h37;
        i_im9 = 8'hAD;
        #10 //22-3
        i_im1 = 8'hAD;
        i_im2 = 8'h3B;
        i_im3 = 8'h3B;
        i_im4 = 8'hBA;
        i_im5 = 8'hB9;
        i_im6 = 8'h39;
        i_im7 = 8'h37;
        i_im8 = 8'hAD;
        i_im9 = 8'h3B;
        #10 //22-4
        i_im1 = 8'h3B;
        i_im2 = 8'h3B;
        i_im3 = 8'h39;
        i_im4 = 8'hB9;
        i_im5 = 8'h39;
        i_im6 = 8'h38;
        i_im7 = 8'hAD;
        i_im8 = 8'h3B;
        i_im9 = 8'hBA;
        #10 //22-5
        i_im1 = 8'h3B;
        i_im2 = 8'h39;
        i_im3 = 8'h37;
        i_im4 = 8'h39;
        i_im5 = 8'h38;
        i_im6 = 8'hB5;
        i_im7 = 8'h3B;
        i_im8 = 8'hBA;
        i_im9 = 8'h2B;
        #10 //22-6
        i_im1 = 8'h39;
        i_im2 = 8'h37;
        i_im3 = 8'h3B;
        i_im4 = 8'h38;
        i_im5 = 8'hB5;
        i_im6 = 8'hB6;
        i_im7 = 8'hBA;
        i_im8 = 8'h2B;
        i_im9 = 8'hB8;
        #10 //22-7
        i_im1 = 8'h37;
        i_im2 = 8'h3B;
        i_im3 = 8'hB8;
        i_im4 = 8'hB5;
        i_im5 = 8'hB6;
        i_im6 = 8'hBB;
        i_im7 = 8'h2B;
        i_im8 = 8'hB8;
        i_im9 = 8'hB7;
        #10 //22-8
        i_im1 = 8'h3B;
        i_im2 = 8'hB8;
        i_im3 = 8'h39;
        i_im4 = 8'hB6;
        i_im5 = 8'hBB;
        i_im6 = 8'h3B;
        i_im7 = 8'hB8;
        i_im8 = 8'hB7;
        i_im9 = 8'h3B;
        #10 //22-9
        i_im1 = 8'hB8;
        i_im2 = 8'h39;
        i_im3 = 8'hB6;
        i_im4 = 8'hBB;
        i_im5 = 8'h3B;
        i_im6 = 8'h39;
        i_im7 = 8'hB7;
        i_im8 = 8'h3B;
        i_im9 = 8'hBC;
        #10 //22-10
        i_im1 = 8'h39;
        i_im2 = 8'hB6;
        i_im3 = 8'hB6;
        i_im4 = 8'h3B;
        i_im5 = 8'h39;
        i_im6 = 8'h3B;
        i_im7 = 8'h3B;
        i_im8 = 8'hBC;
        i_im9 = 8'hAE;
        #10 //22-11
        i_im1 = 8'hB6;
        i_im2 = 8'hB6;
        i_im3 = 8'hA0;
        i_im4 = 8'h39;
        i_im5 = 8'h3B;
        i_im6 = 8'hB0;
        i_im7 = 8'hBC;
        i_im8 = 8'hAE;
        i_im9 = 8'h3B;
        #10 //22-12
        i_im1 = 8'hB6;
        i_im2 = 8'hA0;
        i_im3 = 8'h38;
        i_im4 = 8'h3B;
        i_im5 = 8'hB0;
        i_im6 = 8'hBC;
        i_im7 = 8'hAE;
        i_im8 = 8'h3B;
        i_im9 = 8'h29;
        #10 //22-13
        i_im1 = 8'hA0;
        i_im2 = 8'h38;
        i_im3 = 8'h3B;
        i_im4 = 8'hB0;
        i_im5 = 8'hBC;
        i_im6 = 8'hB5;
        i_im7 = 8'h3B;
        i_im8 = 8'h29;
        i_im9 = 8'hB9;
        #10 //22-14
        i_im1 = 8'h38;
        i_im2 = 8'h3B;
        i_im3 = 8'h38;
        i_im4 = 8'hBC;
        i_im5 = 8'hB5;
        i_im6 = 8'hB4;
        i_im7 = 8'h29;
        i_im8 = 8'hB9;
        i_im9 = 8'h37;
        #10 //22-15
        i_im1 = 8'h3B;
        i_im2 = 8'h38;
        i_im3 = 8'hBB;
        i_im4 = 8'hB5;
        i_im5 = 8'hB4;
        i_im6 = 8'hB9;
        i_im7 = 8'hB9;
        i_im8 = 8'h37;
        i_im9 = 8'h3B;
        #10 //22-16
        i_im1 = 8'h38;
        i_im2 = 8'hBB;
        i_im3 = 8'h39;
        i_im4 = 8'hB4;
        i_im5 = 8'hB9;
        i_im6 = 8'h30;
        i_im7 = 8'h37;
        i_im8 = 8'h3B;
        i_im9 = 8'h34;
        #10 //22-17
        i_im1 = 8'hBB;
        i_im2 = 8'h39;
        i_im3 = 8'h35;
        i_im4 = 8'hB9;
        i_im5 = 8'h30;
        i_im6 = 8'hBA;
        i_im7 = 8'h3B;
        i_im8 = 8'h34;
        i_im9 = 8'hB6;
        #10 //22-18
        i_im1 = 8'h39;
        i_im2 = 8'h35;
        i_im3 = 8'hAF;
        i_im4 = 8'h30;
        i_im5 = 8'hBA;
        i_im6 = 8'h39;
        i_im7 = 8'h34;
        i_im8 = 8'hB6;
        i_im9 = 8'h36;
        #10 //22-19
        i_im1 = 8'h35;
        i_im2 = 8'hAF;
        i_im3 = 8'hB8;
        i_im4 = 8'hBA;
        i_im5 = 8'h39;
        i_im6 = 8'hB8;
        i_im7 = 8'hB6;
        i_im8 = 8'h36;
        i_im9 = 8'h3B;
        #10 //22-20
        i_im1 = 8'hAF;
        i_im2 = 8'hB8;
        i_im3 = 8'h38;
        i_im4 = 8'h39;
        i_im5 = 8'hB8;
        i_im6 = 8'hBB;
        i_im7 = 8'h36;
        i_im8 = 8'h3B;
        i_im9 = 8'h38;
        #10 //22-21
        i_im1 = 8'hB8;
        i_im2 = 8'h38;
        i_im3 = 8'h3A;
        i_im4 = 8'hB8;
        i_im5 = 8'hBB;
        i_im6 = 8'h3B;
        i_im7 = 8'h3B;
        i_im8 = 8'h38;
        i_im9 = 8'hB3;
        #10 //22-22
        i_im1 = 8'h38;
        i_im2 = 8'h3A;
        i_im3 = 8'h38;
        i_im4 = 8'hBB;
        i_im5 = 8'h3B;
        i_im6 = 8'h35;
        i_im7 = 8'h38;
        i_im8 = 8'hB3;
        i_im9 = 8'hB1;
        #10 //22-23
        i_im1 = 8'h3A;
        i_im2 = 8'h38;
        i_im3 = 8'hAE;
        i_im4 = 8'h3B;
        i_im5 = 8'h35;
        i_im6 = 8'h3C;
        i_im7 = 8'hB3;
        i_im8 = 8'hB1;
        i_im9 = 8'hB1;
        #10 //22-24
        i_im1 = 8'h38;
        i_im2 = 8'hAE;
        i_im3 = 8'h34;
        i_im4 = 8'h35;
        i_im5 = 8'h3C;
        i_im6 = 8'h39;
        i_im7 = 8'hB1;
        i_im8 = 8'hB1;
        i_im9 = 8'hB4;
        #10 //22-25
        i_im1 = 8'hAE;
        i_im2 = 8'h34;
        i_im3 = 8'h36;
        i_im4 = 8'h3C;
        i_im5 = 8'h39;
        i_im6 = 8'h3A;
        i_im7 = 8'hB1;
        i_im8 = 8'hB4;
        i_im9 = 8'h2E;
        #10 //22-26
        i_im1 = 8'h34;
        i_im2 = 8'h36;
        i_im3 = 8'h39;
        i_im4 = 8'h39;
        i_im5 = 8'h3A;
        i_im6 = 8'hB2;
        i_im7 = 8'hB4;
        i_im8 = 8'h2E;
        i_im9 = 8'h37;
        #10 //23-1
        i_im1 = 8'h39;
        i_im2 = 8'hB6;
        i_im3 = 8'hBA;
        i_im4 = 8'hBA;
        i_im5 = 8'h36;
        i_im6 = 8'h37;
        i_im7 = 8'h37;
        i_im8 = 8'hAA;
        i_im9 = 8'h39;
        #10 //23-2
        i_im1 = 8'hB6;
        i_im2 = 8'hBA;
        i_im3 = 8'hB9;
        i_im4 = 8'h36;
        i_im5 = 8'h37;
        i_im6 = 8'hAD;
        i_im7 = 8'hAA;
        i_im8 = 8'h39;
        i_im9 = 8'hBA;
        #10 //23-3
        i_im1 = 8'hBA;
        i_im2 = 8'hB9;
        i_im3 = 8'h39;
        i_im4 = 8'h37;
        i_im5 = 8'hAD;
        i_im6 = 8'h3B;
        i_im7 = 8'h39;
        i_im8 = 8'hBA;
        i_im9 = 8'h3B;
        #10 //23-4
        i_im1 = 8'hB9;
        i_im2 = 8'h39;
        i_im3 = 8'h38;
        i_im4 = 8'hAD;
        i_im5 = 8'h3B;
        i_im6 = 8'hBA;
        i_im7 = 8'hBA;
        i_im8 = 8'h3B;
        i_im9 = 8'h3C;
        #10 //23-5
        i_im1 = 8'h39;
        i_im2 = 8'h38;
        i_im3 = 8'hB5;
        i_im4 = 8'h3B;
        i_im5 = 8'hBA;
        i_im6 = 8'h2B;
        i_im7 = 8'h3B;
        i_im8 = 8'h3C;
        i_im9 = 8'hB5;
        #10 //23-6
        i_im1 = 8'h38;
        i_im2 = 8'hB5;
        i_im3 = 8'hB6;
        i_im4 = 8'hBA;
        i_im5 = 8'h2B;
        i_im6 = 8'hB8;
        i_im7 = 8'h3C;
        i_im8 = 8'hB5;
        i_im9 = 8'hB8;
        #10 //23-7
        i_im1 = 8'hB5;
        i_im2 = 8'hB6;
        i_im3 = 8'hBB;
        i_im4 = 8'h2B;
        i_im5 = 8'hB8;
        i_im6 = 8'hB7;
        i_im7 = 8'hB5;
        i_im8 = 8'hB8;
        i_im9 = 8'hB1;
        #10 //23-8
        i_im1 = 8'hB6;
        i_im2 = 8'hBB;
        i_im3 = 8'h3B;
        i_im4 = 8'hB8;
        i_im5 = 8'hB7;
        i_im6 = 8'h3B;
        i_im7 = 8'hB8;
        i_im8 = 8'hB1;
        i_im9 = 8'hA8;
        #10 //23-9
        i_im1 = 8'hBB;
        i_im2 = 8'h3B;
        i_im3 = 8'h39;
        i_im4 = 8'hB7;
        i_im5 = 8'h3B;
        i_im6 = 8'hBC;
        i_im7 = 8'hB1;
        i_im8 = 8'hA8;
        i_im9 = 8'h2F;
        #10 //23-10
        i_im1 = 8'h3B;
        i_im2 = 8'h39;
        i_im3 = 8'h3B;
        i_im4 = 8'h3B;
        i_im5 = 8'hBC;
        i_im6 = 8'hAE;
        i_im7 = 8'hA8;
        i_im8 = 8'h2F;
        i_im9 = 8'h35;
        #10 //23-11
        i_im1 = 8'h39;
        i_im2 = 8'h3B;
        i_im3 = 8'hB0;
        i_im4 = 8'hBC;
        i_im5 = 8'hAE;
        i_im6 = 8'h3B;
        i_im7 = 8'h2F;
        i_im8 = 8'h35;
        i_im9 = 8'hB5;
        #10 //23-12
        i_im1 = 8'h3B;
        i_im2 = 8'hB0;
        i_im3 = 8'hBC;
        i_im4 = 8'hAE;
        i_im5 = 8'h3B;
        i_im6 = 8'h29;
        i_im7 = 8'h35;
        i_im8 = 8'hB5;
        i_im9 = 8'hB4;
        #10 //23-13
        i_im1 = 8'hB0;
        i_im2 = 8'hBC;
        i_im3 = 8'hB5;
        i_im4 = 8'h3B;
        i_im5 = 8'h29;
        i_im6 = 8'hB9;
        i_im7 = 8'hB5;
        i_im8 = 8'hB4;
        i_im9 = 8'hB0;
        #10 //23-14
        i_im1 = 8'hBC;
        i_im2 = 8'hB5;
        i_im3 = 8'hB4;
        i_im4 = 8'h29;
        i_im5 = 8'hB9;
        i_im6 = 8'h37;
        i_im7 = 8'hB4;
        i_im8 = 8'hB0;
        i_im9 = 8'hBA;
        #10 //23-15
        i_im1 = 8'hB5;
        i_im2 = 8'hB4;
        i_im3 = 8'hB9;
        i_im4 = 8'hB9;
        i_im5 = 8'h37;
        i_im6 = 8'h3B;
        i_im7 = 8'hB0;
        i_im8 = 8'hBA;
        i_im9 = 8'h37;
        #10 //23-16
        i_im1 = 8'hB4;
        i_im2 = 8'hB9;
        i_im3 = 8'h30;
        i_im4 = 8'h37;
        i_im5 = 8'h3B;
        i_im6 = 8'h34;
        i_im7 = 8'hBA;
        i_im8 = 8'h37;
        i_im9 = 8'hBA;
        #10 //23-17
        i_im1 = 8'hB9;
        i_im2 = 8'h30;
        i_im3 = 8'hBA;
        i_im4 = 8'h3B;
        i_im5 = 8'h34;
        i_im6 = 8'hB6;
        i_im7 = 8'h37;
        i_im8 = 8'hBA;
        i_im9 = 8'h3B;
        #10 //23-18
        i_im1 = 8'h30;
        i_im2 = 8'hBA;
        i_im3 = 8'h39;
        i_im4 = 8'h34;
        i_im5 = 8'hB6;
        i_im6 = 8'h36;
        i_im7 = 8'hBA;
        i_im8 = 8'h3B;
        i_im9 = 8'h39;
        #10 //23-19
        i_im1 = 8'hBA;
        i_im2 = 8'h39;
        i_im3 = 8'hB8;
        i_im4 = 8'hB6;
        i_im5 = 8'h36;
        i_im6 = 8'h3B;
        i_im7 = 8'h3B;
        i_im8 = 8'h39;
        i_im9 = 8'hB7;
        #10 //23-20
        i_im1 = 8'h39;
        i_im2 = 8'hB8;
        i_im3 = 8'hBB;
        i_im4 = 8'h36;
        i_im5 = 8'h3B;
        i_im6 = 8'h38;
        i_im7 = 8'h39;
        i_im8 = 8'hB7;
        i_im9 = 8'hB9;
        #10 //23-21
        i_im1 = 8'hB8;
        i_im2 = 8'hBB;
        i_im3 = 8'h3B;
        i_im4 = 8'h3B;
        i_im5 = 8'h38;
        i_im6 = 8'hB3;
        i_im7 = 8'hB7;
        i_im8 = 8'hB9;
        i_im9 = 8'h3C;
        #10 //23-22
        i_im1 = 8'hBB;
        i_im2 = 8'h3B;
        i_im3 = 8'h35;
        i_im4 = 8'h38;
        i_im5 = 8'hB3;
        i_im6 = 8'hB1;
        i_im7 = 8'hB9;
        i_im8 = 8'h3C;
        i_im9 = 8'h39;
        #10 //23-23
        i_im1 = 8'h3B;
        i_im2 = 8'h35;
        i_im3 = 8'h3C;
        i_im4 = 8'hB3;
        i_im5 = 8'hB1;
        i_im6 = 8'hB1;
        i_im7 = 8'h3C;
        i_im8 = 8'h39;
        i_im9 = 8'hB9;
        #10 //23-24
        i_im1 = 8'h35;
        i_im2 = 8'h3C;
        i_im3 = 8'h39;
        i_im4 = 8'hB1;
        i_im5 = 8'hB1;
        i_im6 = 8'hB4;
        i_im7 = 8'h39;
        i_im8 = 8'hB9;
        i_im9 = 8'h3B;
        #10 //23-25
        i_im1 = 8'h3C;
        i_im2 = 8'h39;
        i_im3 = 8'h3A;
        i_im4 = 8'hB1;
        i_im5 = 8'hB4;
        i_im6 = 8'h2E;
        i_im7 = 8'hB9;
        i_im8 = 8'h3B;
        i_im9 = 8'h39;
        #10 //23-26
        i_im1 = 8'h39;
        i_im2 = 8'h3A;
        i_im3 = 8'hB2;
        i_im4 = 8'hB4;
        i_im5 = 8'h2E;
        i_im6 = 8'h37;
        i_im7 = 8'h3B;
        i_im8 = 8'h39;
        i_im9 = 8'h36;
        #10 //24-1
        i_im1 = 8'hBA;
        i_im2 = 8'h36;
        i_im3 = 8'h37;
        i_im4 = 8'h37;
        i_im5 = 8'hAA;
        i_im6 = 8'h39;
        i_im7 = 8'hB8;
        i_im8 = 8'h38;
        i_im9 = 8'h39;
        #10 //24-2
        i_im1 = 8'h36;
        i_im2 = 8'h37;
        i_im3 = 8'hAD;
        i_im4 = 8'hAA;
        i_im5 = 8'h39;
        i_im6 = 8'hBA;
        i_im7 = 8'h38;
        i_im8 = 8'h39;
        i_im9 = 8'h39;
        #10 //24-3
        i_im1 = 8'h37;
        i_im2 = 8'hAD;
        i_im3 = 8'h3B;
        i_im4 = 8'h39;
        i_im5 = 8'hBA;
        i_im6 = 8'h3B;
        i_im7 = 8'h39;
        i_im8 = 8'h39;
        i_im9 = 8'hB8;
        #10 //24-4
        i_im1 = 8'hAD;
        i_im2 = 8'h3B;
        i_im3 = 8'hBA;
        i_im4 = 8'hBA;
        i_im5 = 8'h3B;
        i_im6 = 8'h3C;
        i_im7 = 8'h39;
        i_im8 = 8'hB8;
        i_im9 = 8'h3A;
        #10 //24-5
        i_im1 = 8'h3B;
        i_im2 = 8'hBA;
        i_im3 = 8'h2B;
        i_im4 = 8'h3B;
        i_im5 = 8'h3C;
        i_im6 = 8'hB5;
        i_im7 = 8'hB8;
        i_im8 = 8'h3A;
        i_im9 = 8'hBB;
        #10 //24-6
        i_im1 = 8'hBA;
        i_im2 = 8'h2B;
        i_im3 = 8'hB8;
        i_im4 = 8'h3C;
        i_im5 = 8'hB5;
        i_im6 = 8'hB8;
        i_im7 = 8'h3A;
        i_im8 = 8'hBB;
        i_im9 = 8'hBC;
        #10 //24-7
        i_im1 = 8'h2B;
        i_im2 = 8'hB8;
        i_im3 = 8'hB7;
        i_im4 = 8'hB5;
        i_im5 = 8'hB8;
        i_im6 = 8'hB1;
        i_im7 = 8'hBB;
        i_im8 = 8'hBC;
        i_im9 = 8'hB9;
        #10 //24-8
        i_im1 = 8'hB8;
        i_im2 = 8'hB7;
        i_im3 = 8'h3B;
        i_im4 = 8'hB8;
        i_im5 = 8'hB1;
        i_im6 = 8'hA8;
        i_im7 = 8'hBC;
        i_im8 = 8'hB9;
        i_im9 = 8'h31;
        #10 //24-9
        i_im1 = 8'hB7;
        i_im2 = 8'h3B;
        i_im3 = 8'hBC;
        i_im4 = 8'hB1;
        i_im5 = 8'hA8;
        i_im6 = 8'h2F;
        i_im7 = 8'hB9;
        i_im8 = 8'h31;
        i_im9 = 8'hBA;
        #10 //24-10
        i_im1 = 8'h3B;
        i_im2 = 8'hBC;
        i_im3 = 8'hAE;
        i_im4 = 8'hA8;
        i_im5 = 8'h2F;
        i_im6 = 8'h35;
        i_im7 = 8'h31;
        i_im8 = 8'hBA;
        i_im9 = 8'hB6;
        #10 //24-11
        i_im1 = 8'hBC;
        i_im2 = 8'hAE;
        i_im3 = 8'h3B;
        i_im4 = 8'h2F;
        i_im5 = 8'h35;
        i_im6 = 8'hB5;
        i_im7 = 8'hBA;
        i_im8 = 8'hB6;
        i_im9 = 8'h34;
        #10 //24-12
        i_im1 = 8'hAE;
        i_im2 = 8'h3B;
        i_im3 = 8'h29;
        i_im4 = 8'h35;
        i_im5 = 8'hB5;
        i_im6 = 8'hB4;
        i_im7 = 8'hB6;
        i_im8 = 8'h34;
        i_im9 = 8'hB9;
        #10 //24-13
        i_im1 = 8'h3B;
        i_im2 = 8'h29;
        i_im3 = 8'hB9;
        i_im4 = 8'hB5;
        i_im5 = 8'hB4;
        i_im6 = 8'hB0;
        i_im7 = 8'h34;
        i_im8 = 8'hB9;
        i_im9 = 8'h3B;
        #10 //24-14
        i_im1 = 8'h29;
        i_im2 = 8'hB9;
        i_im3 = 8'h37;
        i_im4 = 8'hB4;
        i_im5 = 8'hB0;
        i_im6 = 8'hBA;
        i_im7 = 8'hB9;
        i_im8 = 8'h3B;
        i_im9 = 8'h39;
        #10 //24-15
        i_im1 = 8'hB9;
        i_im2 = 8'h37;
        i_im3 = 8'h3B;
        i_im4 = 8'hB0;
        i_im5 = 8'hBA;
        i_im6 = 8'h37;
        i_im7 = 8'h3B;
        i_im8 = 8'h39;
        i_im9 = 8'hB2;
        #10 //24-16
        i_im1 = 8'h37;
        i_im2 = 8'h3B;
        i_im3 = 8'h34;
        i_im4 = 8'hBA;
        i_im5 = 8'h37;
        i_im6 = 8'hBA;
        i_im7 = 8'h39;
        i_im8 = 8'hB2;
        i_im9 = 8'h3A;
        #10 //24-17
        i_im1 = 8'h3B;
        i_im2 = 8'h34;
        i_im3 = 8'hB6;
        i_im4 = 8'h37;
        i_im5 = 8'hBA;
        i_im6 = 8'h3B;
        i_im7 = 8'hB2;
        i_im8 = 8'h3A;
        i_im9 = 8'hBB;
        #10 //24-18
        i_im1 = 8'h34;
        i_im2 = 8'hB6;
        i_im3 = 8'h36;
        i_im4 = 8'hBA;
        i_im5 = 8'h3B;
        i_im6 = 8'h39;
        i_im7 = 8'h3A;
        i_im8 = 8'hBB;
        i_im9 = 8'h2C;
        #10 //24-19
        i_im1 = 8'hB6;
        i_im2 = 8'h36;
        i_im3 = 8'h3B;
        i_im4 = 8'h3B;
        i_im5 = 8'h39;
        i_im6 = 8'hB7;
        i_im7 = 8'hBB;
        i_im8 = 8'h2C;
        i_im9 = 8'hB3;
        #10 //24-20
        i_im1 = 8'h36;
        i_im2 = 8'h3B;
        i_im3 = 8'h38;
        i_im4 = 8'h39;
        i_im5 = 8'hB7;
        i_im6 = 8'hB9;
        i_im7 = 8'h2C;
        i_im8 = 8'hB3;
        i_im9 = 8'hBB;
        #10 //24-21
        i_im1 = 8'h3B;
        i_im2 = 8'h38;
        i_im3 = 8'hB3;
        i_im4 = 8'hB7;
        i_im5 = 8'hB9;
        i_im6 = 8'h3C;
        i_im7 = 8'hB3;
        i_im8 = 8'hBB;
        i_im9 = 8'h3A;
        #10 //24-22
        i_im1 = 8'h38;
        i_im2 = 8'hB3;
        i_im3 = 8'hB1;
        i_im4 = 8'hB9;
        i_im5 = 8'h3C;
        i_im6 = 8'h39;
        i_im7 = 8'hBB;
        i_im8 = 8'h3A;
        i_im9 = 8'h37;
        #10 //24-23
        i_im1 = 8'hB3;
        i_im2 = 8'hB1;
        i_im3 = 8'hB1;
        i_im4 = 8'h3C;
        i_im5 = 8'h39;
        i_im6 = 8'hB9;
        i_im7 = 8'h3A;
        i_im8 = 8'h37;
        i_im9 = 8'h3A;
        #10 //24-24
        i_im1 = 8'hB1;
        i_im2 = 8'hB1;
        i_im3 = 8'hB4;
        i_im4 = 8'h39;
        i_im5 = 8'hB9;
        i_im6 = 8'h3B;
        i_im7 = 8'h37;
        i_im8 = 8'h3A;
        i_im9 = 8'hBC;
        #10 //24-25
        i_im1 = 8'hB1;
        i_im2 = 8'hB4;
        i_im3 = 8'h2E;
        i_im4 = 8'hB9;
        i_im5 = 8'h3B;
        i_im6 = 8'h39;
        i_im7 = 8'h3A;
        i_im8 = 8'hBC;
        i_im9 = 8'h35;
        #10 //24-26
        i_im1 = 8'hB4;
        i_im2 = 8'h2E;
        i_im3 = 8'h37;
        i_im4 = 8'h3B;
        i_im5 = 8'h39;
        i_im6 = 8'h36;
        i_im7 = 8'hBC;
        i_im8 = 8'h35;
        i_im9 = 8'h2C;
        #10 //25-1
        i_im1 = 8'h37;
        i_im2 = 8'hAA;
        i_im3 = 8'h39;
        i_im4 = 8'hB8;
        i_im5 = 8'h38;
        i_im6 = 8'h39;
        i_im7 = 8'h39;
        i_im8 = 8'hB9;
        i_im9 = 8'h36;
        #10 //25-2
        i_im1 = 8'hAA;
        i_im2 = 8'h39;
        i_im3 = 8'hBA;
        i_im4 = 8'h38;
        i_im5 = 8'h39;
        i_im6 = 8'h39;
        i_im7 = 8'hB9;
        i_im8 = 8'h36;
        i_im9 = 8'hBB;
        #10 //25-3
        i_im1 = 8'h39;
        i_im2 = 8'hBA;
        i_im3 = 8'h3B;
        i_im4 = 8'h39;
        i_im5 = 8'h39;
        i_im6 = 8'hB8;
        i_im7 = 8'h36;
        i_im8 = 8'hBB;
        i_im9 = 8'h32;
        #10 //25-4
        i_im1 = 8'hBA;
        i_im2 = 8'h3B;
        i_im3 = 8'h3C;
        i_im4 = 8'h39;
        i_im5 = 8'hB8;
        i_im6 = 8'h3A;
        i_im7 = 8'hBB;
        i_im8 = 8'h32;
        i_im9 = 8'hB7;
        #10 //25-5
        i_im1 = 8'h3B;
        i_im2 = 8'h3C;
        i_im3 = 8'hB5;
        i_im4 = 8'hB8;
        i_im5 = 8'h3A;
        i_im6 = 8'hBB;
        i_im7 = 8'h32;
        i_im8 = 8'hB7;
        i_im9 = 8'h3A;
        #10 //25-6
        i_im1 = 8'h3C;
        i_im2 = 8'hB5;
        i_im3 = 8'hB8;
        i_im4 = 8'h3A;
        i_im5 = 8'hBB;
        i_im6 = 8'hBC;
        i_im7 = 8'hB7;
        i_im8 = 8'h3A;
        i_im9 = 8'h31;
        #10 //25-7
        i_im1 = 8'hB5;
        i_im2 = 8'hB8;
        i_im3 = 8'hB1;
        i_im4 = 8'hBB;
        i_im5 = 8'hBC;
        i_im6 = 8'hB9;
        i_im7 = 8'h3A;
        i_im8 = 8'h31;
        i_im9 = 8'h3C;
        #10 //25-8
        i_im1 = 8'hB8;
        i_im2 = 8'hB1;
        i_im3 = 8'hA8;
        i_im4 = 8'hBC;
        i_im5 = 8'hB9;
        i_im6 = 8'h31;
        i_im7 = 8'h31;
        i_im8 = 8'h3C;
        i_im9 = 8'h32;
        #10 //25-9
        i_im1 = 8'hB1;
        i_im2 = 8'hA8;
        i_im3 = 8'h2F;
        i_im4 = 8'hB9;
        i_im5 = 8'h31;
        i_im6 = 8'hBA;
        i_im7 = 8'h3C;
        i_im8 = 8'h32;
        i_im9 = 8'h3C;
        #10 //25-10
        i_im1 = 8'hA8;
        i_im2 = 8'h2F;
        i_im3 = 8'h35;
        i_im4 = 8'h31;
        i_im5 = 8'hBA;
        i_im6 = 8'hB6;
        i_im7 = 8'h32;
        i_im8 = 8'h3C;
        i_im9 = 8'h39;
        #10 //25-11
        i_im1 = 8'h2F;
        i_im2 = 8'h35;
        i_im3 = 8'hB5;
        i_im4 = 8'hBA;
        i_im5 = 8'hB6;
        i_im6 = 8'h34;
        i_im7 = 8'h3C;
        i_im8 = 8'h39;
        i_im9 = 8'h37;
        #10 //25-12
        i_im1 = 8'h35;
        i_im2 = 8'hB5;
        i_im3 = 8'hB4;
        i_im4 = 8'hB6;
        i_im5 = 8'h34;
        i_im6 = 8'hB9;
        i_im7 = 8'h39;
        i_im8 = 8'h37;
        i_im9 = 8'h3A;
        #10 //25-13
        i_im1 = 8'hB5;
        i_im2 = 8'hB4;
        i_im3 = 8'hB0;
        i_im4 = 8'h34;
        i_im5 = 8'hB9;
        i_im6 = 8'h3B;
        i_im7 = 8'h37;
        i_im8 = 8'h3A;
        i_im9 = 8'h39;
        #10 //25-14
        i_im1 = 8'hB4;
        i_im2 = 8'hB0;
        i_im3 = 8'hBA;
        i_im4 = 8'hB9;
        i_im5 = 8'h3B;
        i_im6 = 8'h39;
        i_im7 = 8'h3A;
        i_im8 = 8'h39;
        i_im9 = 8'h2F;
        #10 //25-15
        i_im1 = 8'hB0;
        i_im2 = 8'hBA;
        i_im3 = 8'h37;
        i_im4 = 8'h3B;
        i_im5 = 8'h39;
        i_im6 = 8'hB2;
        i_im7 = 8'h39;
        i_im8 = 8'h2F;
        i_im9 = 8'hB9;
        #10 //25-16
        i_im1 = 8'hBA;
        i_im2 = 8'h37;
        i_im3 = 8'hBA;
        i_im4 = 8'h39;
        i_im5 = 8'hB2;
        i_im6 = 8'h3A;
        i_im7 = 8'h2F;
        i_im8 = 8'hB9;
        i_im9 = 8'hB8;
        #10 //25-17
        i_im1 = 8'h37;
        i_im2 = 8'hBA;
        i_im3 = 8'h3B;
        i_im4 = 8'hB2;
        i_im5 = 8'h3A;
        i_im6 = 8'hBB;
        i_im7 = 8'hB9;
        i_im8 = 8'hB8;
        i_im9 = 8'hB2;
        #10 //25-18
        i_im1 = 8'hBA;
        i_im2 = 8'h3B;
        i_im3 = 8'h39;
        i_im4 = 8'h3A;
        i_im5 = 8'hBB;
        i_im6 = 8'h2C;
        i_im7 = 8'hB8;
        i_im8 = 8'hB2;
        i_im9 = 8'h39;
        #10 //25-19
        i_im1 = 8'h3B;
        i_im2 = 8'h39;
        i_im3 = 8'hB7;
        i_im4 = 8'hBB;
        i_im5 = 8'h2C;
        i_im6 = 8'hB3;
        i_im7 = 8'hB2;
        i_im8 = 8'h39;
        i_im9 = 8'h29;
        #10 //25-20
        i_im1 = 8'h39;
        i_im2 = 8'hB7;
        i_im3 = 8'hB9;
        i_im4 = 8'h2C;
        i_im5 = 8'hB3;
        i_im6 = 8'hBB;
        i_im7 = 8'h39;
        i_im8 = 8'h29;
        i_im9 = 8'hBA;
        #10 //25-21
        i_im1 = 8'hB7;
        i_im2 = 8'hB9;
        i_im3 = 8'h3C;
        i_im4 = 8'hB3;
        i_im5 = 8'hBB;
        i_im6 = 8'h3A;
        i_im7 = 8'h29;
        i_im8 = 8'hBA;
        i_im9 = 8'h3B;
        #10 //25-22
        i_im1 = 8'hB9;
        i_im2 = 8'h3C;
        i_im3 = 8'h39;
        i_im4 = 8'hBB;
        i_im5 = 8'h3A;
        i_im6 = 8'h37;
        i_im7 = 8'hBA;
        i_im8 = 8'h3B;
        i_im9 = 8'hB9;
        #10 //25-23
        i_im1 = 8'h3C;
        i_im2 = 8'h39;
        i_im3 = 8'hB9;
        i_im4 = 8'h3A;
        i_im5 = 8'h37;
        i_im6 = 8'h3A;
        i_im7 = 8'h3B;
        i_im8 = 8'hB9;
        i_im9 = 8'hB5;
        #10 //25-24
        i_im1 = 8'h39;
        i_im2 = 8'hB9;
        i_im3 = 8'h3B;
        i_im4 = 8'h37;
        i_im5 = 8'h3A;
        i_im6 = 8'hBC;
        i_im7 = 8'hB9;
        i_im8 = 8'hB5;
        i_im9 = 8'hBA;
        #10 //25-25
        i_im1 = 8'hB9;
        i_im2 = 8'h3B;
        i_im3 = 8'h39;
        i_im4 = 8'h3A;
        i_im5 = 8'hBC;
        i_im6 = 8'h35;
        i_im7 = 8'hB5;
        i_im8 = 8'hBA;
        i_im9 = 8'h3A;
        #10 //25-26
        i_im1 = 8'h3B;
        i_im2 = 8'h39;
        i_im3 = 8'h36;
        i_im4 = 8'hBC;
        i_im5 = 8'h35;
        i_im6 = 8'h2C;
        i_im7 = 8'hBA;
        i_im8 = 8'h3A;
        i_im9 = 8'hB7;
        #10 //26-1
        i_im1 = 8'hB8;
        i_im2 = 8'h38;
        i_im3 = 8'h39;
        i_im4 = 8'h39;
        i_im5 = 8'hB9;
        i_im6 = 8'h36;
        i_im7 = 8'h37;
        i_im8 = 8'h25;
        i_im9 = 8'h2A;
        #10 //26-2
        i_im1 = 8'h38;
        i_im2 = 8'h39;
        i_im3 = 8'h39;
        i_im4 = 8'hB9;
        i_im5 = 8'h36;
        i_im6 = 8'hBB;
        i_im7 = 8'h25;
        i_im8 = 8'h2A;
        i_im9 = 8'h3A;
        #10 //26-3
        i_im1 = 8'h39;
        i_im2 = 8'h39;
        i_im3 = 8'hB8;
        i_im4 = 8'h36;
        i_im5 = 8'hBB;
        i_im6 = 8'h32;
        i_im7 = 8'h2A;
        i_im8 = 8'h3A;
        i_im9 = 8'h3B;
        #10 //26-4
        i_im1 = 8'h39;
        i_im2 = 8'hB8;
        i_im3 = 8'h3A;
        i_im4 = 8'hBB;
        i_im5 = 8'h32;
        i_im6 = 8'hB7;
        i_im7 = 8'h3A;
        i_im8 = 8'h3B;
        i_im9 = 8'hB7;
        #10 //26-5
        i_im1 = 8'hB8;
        i_im2 = 8'h3A;
        i_im3 = 8'hBB;
        i_im4 = 8'h32;
        i_im5 = 8'hB7;
        i_im6 = 8'h3A;
        i_im7 = 8'h3B;
        i_im8 = 8'hB7;
        i_im9 = 8'hBA;
        #10 //26-6
        i_im1 = 8'h3A;
        i_im2 = 8'hBB;
        i_im3 = 8'hBC;
        i_im4 = 8'hB7;
        i_im5 = 8'h3A;
        i_im6 = 8'h31;
        i_im7 = 8'hB7;
        i_im8 = 8'hBA;
        i_im9 = 8'hB9;
        #10 //26-7
        i_im1 = 8'hBB;
        i_im2 = 8'hBC;
        i_im3 = 8'hB9;
        i_im4 = 8'h3A;
        i_im5 = 8'h31;
        i_im6 = 8'h3C;
        i_im7 = 8'hBA;
        i_im8 = 8'hB9;
        i_im9 = 8'h2E;
        #10 //26-8
        i_im1 = 8'hBC;
        i_im2 = 8'hB9;
        i_im3 = 8'h31;
        i_im4 = 8'h31;
        i_im5 = 8'h3C;
        i_im6 = 8'h32;
        i_im7 = 8'hB9;
        i_im8 = 8'h2E;
        i_im9 = 8'h3B;
        #10 //26-9
        i_im1 = 8'hB9;
        i_im2 = 8'h31;
        i_im3 = 8'hBA;
        i_im4 = 8'h3C;
        i_im5 = 8'h32;
        i_im6 = 8'h3C;
        i_im7 = 8'h2E;
        i_im8 = 8'h3B;
        i_im9 = 8'hBB;
        #10 //26-10
        i_im1 = 8'h31;
        i_im2 = 8'hBA;
        i_im3 = 8'hB6;
        i_im4 = 8'h32;
        i_im5 = 8'h3C;
        i_im6 = 8'h39;
        i_im7 = 8'h3B;
        i_im8 = 8'hBB;
        i_im9 = 8'hBC;
        #10 //26-11
        i_im1 = 8'hBA;
        i_im2 = 8'hB6;
        i_im3 = 8'h34;
        i_im4 = 8'h3C;
        i_im5 = 8'h39;
        i_im6 = 8'h37;
        i_im7 = 8'hBB;
        i_im8 = 8'hBC;
        i_im9 = 8'hB7;
        #10 //26-12
        i_im1 = 8'hB6;
        i_im2 = 8'h34;
        i_im3 = 8'hB9;
        i_im4 = 8'h39;
        i_im5 = 8'h37;
        i_im6 = 8'h3A;
        i_im7 = 8'hBC;
        i_im8 = 8'hB7;
        i_im9 = 8'h3A;
        #10 //26-13
        i_im1 = 8'h34;
        i_im2 = 8'hB9;
        i_im3 = 8'h3B;
        i_im4 = 8'h37;
        i_im5 = 8'h3A;
        i_im6 = 8'h39;
        i_im7 = 8'hB7;
        i_im8 = 8'h3A;
        i_im9 = 8'h3B;
        #10 //26-14
        i_im1 = 8'hB9;
        i_im2 = 8'h3B;
        i_im3 = 8'h39;
        i_im4 = 8'h3A;
        i_im5 = 8'h39;
        i_im6 = 8'h2F;
        i_im7 = 8'h3A;
        i_im8 = 8'h3B;
        i_im9 = 8'hB9;
        #10 //26-15
        i_im1 = 8'h3B;
        i_im2 = 8'h39;
        i_im3 = 8'hB2;
        i_im4 = 8'h39;
        i_im5 = 8'h2F;
        i_im6 = 8'hB9;
        i_im7 = 8'h3B;
        i_im8 = 8'hB9;
        i_im9 = 8'hB7;
        #10 //26-16
        i_im1 = 8'h39;
        i_im2 = 8'hB2;
        i_im3 = 8'h3A;
        i_im4 = 8'h2F;
        i_im5 = 8'hB9;
        i_im6 = 8'hB8;
        i_im7 = 8'hB9;
        i_im8 = 8'hB7;
        i_im9 = 8'h00;
        #10 //26-17
        i_im1 = 8'hB2;
        i_im2 = 8'h3A;
        i_im3 = 8'hBB;
        i_im4 = 8'hB9;
        i_im5 = 8'hB8;
        i_im6 = 8'hB2;
        i_im7 = 8'hB7;
        i_im8 = 8'h00;
        i_im9 = 8'hB7;
        #10 //26-18
        i_im1 = 8'h3A;
        i_im2 = 8'hBB;
        i_im3 = 8'h2C;
        i_im4 = 8'hB8;
        i_im5 = 8'hB2;
        i_im6 = 8'h39;
        i_im7 = 8'h00;
        i_im8 = 8'hB7;
        i_im9 = 8'h39;
        #10 //26-19
        i_im1 = 8'hBB;
        i_im2 = 8'h2C;
        i_im3 = 8'hB3;
        i_im4 = 8'hB2;
        i_im5 = 8'h39;
        i_im6 = 8'h29;
        i_im7 = 8'hB7;
        i_im8 = 8'h39;
        i_im9 = 8'hB4;
        #10 //26-20
        i_im1 = 8'h2C;
        i_im2 = 8'hB3;
        i_im3 = 8'hBB;
        i_im4 = 8'h39;
        i_im5 = 8'h29;
        i_im6 = 8'hBA;
        i_im7 = 8'h39;
        i_im8 = 8'hB4;
        i_im9 = 8'hBA;
        #10 //26-21
        i_im1 = 8'hB3;
        i_im2 = 8'hBB;
        i_im3 = 8'h3A;
        i_im4 = 8'h29;
        i_im5 = 8'hBA;
        i_im6 = 8'h3B;
        i_im7 = 8'hB4;
        i_im8 = 8'hBA;
        i_im9 = 8'h37;
        #10 //26-22
        i_im1 = 8'hBB;
        i_im2 = 8'h3A;
        i_im3 = 8'h37;
        i_im4 = 8'hBA;
        i_im5 = 8'h3B;
        i_im6 = 8'hB9;
        i_im7 = 8'hBA;
        i_im8 = 8'h37;
        i_im9 = 8'h39;
        #10 //26-23
        i_im1 = 8'h3A;
        i_im2 = 8'h37;
        i_im3 = 8'h3A;
        i_im4 = 8'h3B;
        i_im5 = 8'hB9;
        i_im6 = 8'hB5;
        i_im7 = 8'h37;
        i_im8 = 8'h39;
        i_im9 = 8'h39;
        #10 //26-24
        i_im1 = 8'h37;
        i_im2 = 8'h3A;
        i_im3 = 8'hBC;
        i_im4 = 8'hB9;
        i_im5 = 8'hB5;
        i_im6 = 8'hBA;
        i_im7 = 8'h39;
        i_im8 = 8'h39;
        i_im9 = 8'hBB;
        #10 //26-25
        i_im1 = 8'h3A;
        i_im2 = 8'hBC;
        i_im3 = 8'h35;
        i_im4 = 8'hB5;
        i_im5 = 8'hBA;
        i_im6 = 8'h3A;
        i_im7 = 8'h39;
        i_im8 = 8'hBB;
        i_im9 = 8'hBC;
        #10 //26-26
        i_im1 = 8'hBC;
        i_im2 = 8'h35;
        i_im3 = 8'h2C;
        i_im4 = 8'hBA;
        i_im5 = 8'h3A;
        i_im6 = 8'hB7;
        i_im7 = 8'hBB;
        i_im8 = 8'hBC;
        i_im9 = 8'h3A;



        #1000 $finish;
    end
    
    always begin
        #5 clk=~clk;
    end

    reg [6:0] count,count_next;
    reg [6:0] row_count,row_count_next;
    always @(*) begin
        row_count_next = row_count;
        if(o_valid) begin
            if(count<=25) begin
                count_next = count+1;
            end
            else begin
                count_next = 1;
                row_count_next = row_count + 1;
            end
        end
        else begin
            count_next = count;
        end
    end
    always @(posedge clk or negedge i_rst_n) begin
        if(!i_rst_n) begin
            count <= 1;
            row_count <= 1;
        end
        else begin
            count <= count_next;
            row_count <= row_count_next;
        end
        
    end

    mac        DUT(.clk(clk),
               .i_rst_n(i_rst_n),
               .i_inhibit(1'b0),
               .i_valid(i_valid),
               .i_q(9'd0),
               .zero_vector(9'd0),

               // input pixels
               .i_im1(i_im1),
               .i_im2(i_im2),
               .i_im3(i_im3),
               .i_im4(i_im4),
               .i_im5(i_im5),
               .i_im6(i_im6),
               .i_im7(i_im7),
               .i_im8(i_im8),
               .i_im9(i_im9),

               // input weights
               .i_ker1(i_ker1),
               .i_ker2(i_ker2),
               .i_ker3(i_ker3),
               .i_ker4(i_ker4),
               .i_ker5(i_ker5),
               .i_ker6(i_ker6),
               .i_ker7(i_ker7),
               .i_ker8(i_ker8),
               .i_ker9(i_ker9),

               // output ports
               .o_valid(o_valid),
               .o_conv(o_conv)
              );
endmodule