module top_module (
    input clk,
    input [7:0] in,
    output [7:0] pedge
);






endmodule
